module font_rom (
    input  wire clk_in, 
    input  wire [8:0] addr,  // 9-bit address for up to 320 rows
    output reg [15:0] data   // 16-bit data output (one row of 16 bits)
);

    logic [15:0] memory [0:319]; // 320 rows of 16-bit data (20 blocks × 16 rows each)

    initial begin
        // Font for 'A' (Block 0, 16×16 grid)
        memory[0]  = 16'b0000011111100000; 
        memory[1]  = 16'b0000110000110000; 
        memory[2]  = 16'b0001100000011000;
        memory[3]  = 16'b0011000000001100;
        memory[4]  = 16'b0011000000001100;
        memory[5]  = 16'b0110000000000110;
        memory[6]  = 16'b0111111111111110; 
        memory[7]  = 16'b1100000000000011; 
        memory[8]  = 16'b1100000000000011;
        memory[9]  = 16'b1100000000000011;
        memory[10] = 16'b1100000000000011;
        memory[11] = 16'b1100000000000011;
        memory[12] = 16'b1100000000000011;
        memory[13] = 16'b1100000000000011;
        memory[14] = 16'b0000000000000000;
        memory[15] = 16'b0000000000000000;

        // Font for 'B' (Block 1, 16×16 grid)
        memory[16] = 16'b1111111111110000;
        memory[17] = 16'b1000000000001000;
        memory[18] = 16'b1000000000000100;
        memory[19] = 16'b1000000000000100;
        memory[20] = 16'b1000000000000100;
        memory[21] = 16'b1000000000001000;
        memory[22] = 16'b1111111111110000;
        memory[23] = 16'b1000000000000100;
        memory[24] = 16'b1000000000000010;
        memory[25] = 16'b1000000000000010;
        memory[26] = 16'b1000000000000010;
        memory[27] = 16'b1000000000000100;
        memory[28] = 16'b1000000000001000;
        memory[29] = 16'b1111111111110000;
        memory[30] = 16'b0000000000000000;
        memory[31] = 16'b0000000000000000;

        //C
        memory[32] = 16'b0000111111111000;
        memory[33] = 16'b0011000000001100;
        memory[34] = 16'b0100000000000010;
        memory[35] = 16'b1000000000000000;
        memory[36] = 16'b1000000000000000;
        memory[37] = 16'b1000000000000000;
        memory[38] = 16'b1000000000000000;
        memory[39] = 16'b1000000000000000;
        memory[40] = 16'b1000000000000000;
        memory[41] = 16'b1000000000000000;
        memory[42] = 16'b1000000000000000;
        memory[43] = 16'b1000000000000000;
        memory[44] = 16'b0100000000000010;
        memory[45] = 16'b0011000000001100;
        memory[46] = 16'b0000111111111000;
        memory[47] = 16'b0000000000000000;

        //D
        memory[48] = 16'b1111111111110000;
        memory[49] = 16'b1000000000001000;
        memory[50] = 16'b1000000000000100;
        memory[51] = 16'b1000000000000010;
        memory[52] = 16'b1000000000000010;
        memory[53] = 16'b1000000000000010;
        memory[54] = 16'b1000000000000010;
        memory[55] = 16'b1000000000000010;
        memory[56] = 16'b1000000000000010;
        memory[57] = 16'b1000000000000010;
        memory[58] = 16'b1000000000000010;
        memory[59] = 16'b1000000000000010;
        memory[60] = 16'b1000000000000100;
        memory[61] = 16'b1000000000001000;
        memory[62] = 16'b1111111111110000;
        memory[63] = 16'b0000000000000000;

        //E
        memory[64] = 16'b1111111111111110;
        memory[65] = 16'b1000000000000000;
        memory[66] = 16'b1000000000000000;
        memory[67] = 16'b1000000000000000;
        memory[68] = 16'b1000000000000000;
        memory[69] = 16'b1111111111111000;
        memory[70] = 16'b1000000000000000;
        memory[71] = 16'b1000000000000000;
        memory[72] = 16'b1000000000000000;
        memory[73] = 16'b1000000000000000;
        memory[74] = 16'b1000000000000000;
        memory[75] = 16'b1111111111111110;
        memory[76] = 16'b0000000000000000;
        memory[77] = 16'b0000000000000000;
        memory[78] = 16'b0000000000000000;
        memory[79] = 16'b0000000000000000;

        //F
        memory[80] = 16'b1111111111111110;
        memory[81] = 16'b1000000000000000;
        memory[82] = 16'b1000000000000000;
        memory[83] = 16'b1000000000000000;
        memory[84] = 16'b1000000000000000;
        memory[85] = 16'b1111111111111000;
        memory[86] = 16'b1000000000000000;
        memory[87] = 16'b1000000000000000;
        memory[88] = 16'b1000000000000000;
        memory[89] = 16'b1000000000000000;
        memory[90] = 16'b1000000000000000;
        memory[91] = 16'b1000000000000000;
        memory[92] = 16'b1000000000000000;
        memory[93] = 16'b0000000000000000;
        memory[94] = 16'b0000000000000000;
        memory[95] = 16'b0000000000000000;

        //G
        memory[96] = 16'b0000111111111000;
        memory[97] = 16'b0011000000001100;
        memory[98] = 16'b0100000000000010;
        memory[99] = 16'b1000000000000000;
        memory[100] = 16'b1000000000000000;
        memory[101] = 16'b1000001111111100;
        memory[102] = 16'b1000000000000010;
        memory[103] = 16'b1000000000000010;
        memory[104] = 16'b1000000000000010;
        memory[105] = 16'b1000000000000010;
        memory[106] = 16'b0100000000000010;
        memory[107] = 16'b0011000000001100;
        memory[108] = 16'b0000111111111000;
        memory[109] = 16'b0000000000000000;
        memory[110] = 16'b0000000000000000;
        memory[111] = 16'b0000000000000000;

        //1
        memory[112] = 16'b0000001000000000;
        memory[113] = 16'b0000011000000000;
        memory[114] = 16'b0000111000000000;
        memory[115] = 16'b0000001000000000;
        memory[116] = 16'b0000001000000000;
        memory[117] = 16'b0000001000000000;
        memory[118] = 16'b0000001000000000;
        memory[119] = 16'b0000001000000000;
        memory[120] = 16'b0000001000000000;
        memory[121] = 16'b0000001000000000;
        memory[122] = 16'b0000001000000000;
        memory[123] = 16'b0000111111111100;
        memory[124] = 16'b0000000000000000;
        memory[125] = 16'b0000000000000000;
        memory[126] = 16'b0000000000000000;
        memory[127] = 16'b0000000000000000;

        //2
        memory[128] = 16'b0000111111110000;
        memory[129] = 16'b0011111111111110;
        memory[130] = 16'b0111000000001110;
        memory[131] = 16'b1100000000000110;
        memory[132] = 16'b0000000000000110;
        memory[133] = 16'b0000000000000110;
        memory[134] = 16'b0000000000000110;
        memory[135] = 16'b0000000000011100;
        memory[136] = 16'b0000000000111000;
        memory[137] = 16'b0000000001110000;
        memory[138] = 16'b0000000011100000;
        memory[139] = 16'b0000000111000000;
        memory[140] = 16'b0000011100000000;
        memory[141] = 16'b0001110000000000;
        memory[142] = 16'b1111111111111110;
        memory[143] = 16'b0000000000000000;

        //3
        memory[144] = 16'b0000111111110000;
        memory[145] = 16'b0011000000001100;
        memory[146] = 16'b0100000000000010;
        memory[147] = 16'b1000000000000010;
        memory[148] = 16'b0000000000000010;
        memory[149] = 16'b0000000000001100;
        memory[150] = 16'b0000001111110000;
        memory[151] = 16'b0000000000001100;
        memory[152] = 16'b0000000000000010;
        memory[153] = 16'b0000000000000010;
        memory[154] = 16'b1000000000000010;
        memory[155] = 16'b0100000000000010;
        memory[156] = 16'b0011000000001100;
        memory[157] = 16'b0000111111110000;
        memory[158] = 16'b0000000000000000;
        memory[159] = 16'b0000000000000000;

        //4
        memory[160] = 16'b0000000000010000;
        memory[161] = 16'b0000000000110000;
        memory[162] = 16'b0000000001010000;
        memory[163] = 16'b0000000010010000;
        memory[164] = 16'b0000000100010000;
        memory[165] = 16'b0000001000010000;
        memory[166] = 16'b0000010000010000;
        memory[167] = 16'b0000100000010000;
        memory[168] = 16'b0001000000010000;
        memory[169] = 16'b0011111111111110;
        memory[170] = 16'b0000000000010000;
        memory[171] = 16'b0000000000010000;
        memory[172] = 16'b0000000000010000;
        memory[173] = 16'b0000000000000000;
        memory[174] = 16'b0000000000000000;
        memory[175] = 16'b0000000000000000;

        //5
        memory[176] = 16'b1111111111111110;
        memory[177] = 16'b1000000000000000;
        memory[178] = 16'b1000000000000000;
        memory[179] = 16'b1000000000000000;
        memory[180] = 16'b1111111111110000;
        memory[181] = 16'b0000000000001100;
        memory[182] = 16'b0000000000000010;
        memory[183] = 16'b0000000000000010;
        memory[184] = 16'b0000000000000010;
        memory[185] = 16'b1000000000000010;
        memory[186] = 16'b0100000000000010;
        memory[187] = 16'b0011000000001100;
        memory[188] = 16'b0000111111110000;
        memory[189] = 16'b0000000000000000;
        memory[190] = 16'b0000000000000000;
        memory[191] = 16'b0000000000000000;

        //6
        memory[192] = 16'b0000001111111000;
        memory[193] = 16'b0000110000001100;
        memory[194] = 16'b0001100000000010;
        memory[195] = 16'b0011000000000000;
        memory[196] = 16'b0111111111111000;
        memory[197] = 16'b1100000000001100;
        memory[198] = 16'b1000000000000010;
        memory[199] = 16'b1000000000000010;
        memory[200] = 16'b1000000000000010;
        memory[201] = 16'b1000000000000010;
        memory[202] = 16'b0100000000000010;
        memory[203] = 16'b0011000000001100;
        memory[204] = 16'b0000111111110000;
        memory[205] = 16'b0000000000000000;
        memory[206] = 16'b0000000000000000;
        memory[207] = 16'b0000000000000000;

        //7
        memory[208] = 16'b1111111111111110;
        memory[209] = 16'b0000000000000010;
        memory[210] = 16'b0000000000000100;
        memory[211] = 16'b0000000000001000;
        memory[212] = 16'b0000000000010000;
        memory[213] = 16'b0000000000100000;
        memory[214] = 16'b0000000001000000;
        memory[215] = 16'b0000000010000000;
        memory[216] = 16'b0000000100000000;
        memory[217] = 16'b0000001000000000;
        memory[218] = 16'b0000010000000000;
        memory[219] = 16'b0000100000000000;
        memory[220] = 16'b0001000000000000;
        memory[221] = 16'b0000000000000000;
        memory[222] = 16'b0000000000000000;
        memory[223] = 16'b0000000000000000;

        //8
        memory[224] = 16'b0000111111110000;
        memory[225] = 16'b0011000000001100;
        memory[226] = 16'b0100000000000010;
        memory[227] = 16'b1000000000000010;
        memory[228] = 16'b1000000000000010;
        memory[229] = 16'b0100000000000010;
        memory[230] = 16'b0011000000001100;
        memory[231] = 16'b0000111111110000;
        memory[232] = 16'b0011000000001100;
        memory[233] = 16'b0100000000000010;
        memory[234] = 16'b1000000000000010;
        memory[235] = 16'b1000000000000010;
        memory[236] = 16'b0100000000000010;
        memory[237] = 16'b0011000000001100;
        memory[238] = 16'b0000111111110000;
        memory[239] = 16'b0000000000000000;

        //9
        memory[240] = 16'b0000111111110000;
        memory[241] = 16'b0011000000001100;
        memory[242] = 16'b0100000000000010;
        memory[243] = 16'b1000000000000010;
        memory[244] = 16'b1000000000000010;
        memory[245] = 16'b1000000000000010;
        memory[246] = 16'b0100000000000010;
        memory[247] = 16'b0011111111111110;
        memory[248] = 16'b0000000000000010;
        memory[249] = 16'b0000000000000010;
        memory[250] = 16'b0000000000000010;
        memory[251] = 16'b1000000000000100;
        memory[252] = 16'b0100000000001000;
        memory[253] = 16'b0011000000110000;
        memory[254] = 16'b0000111111000000;
        memory[255] = 16'b0000000000000000;

        //blank
        // Blank sprite starting at address 256
        memory[256] = 16'b0000000000000000;
        memory[257] = 16'b0000000000000000;
        memory[258] = 16'b0000000000000000;
        memory[259] = 16'b0000000000000000;
        memory[260] = 16'b0000000000000000;
        memory[261] = 16'b0000000000000000;
        memory[262] = 16'b0000000000000000;
        memory[263] = 16'b0000000000000000;
        memory[264] = 16'b0000000000000000;
        memory[265] = 16'b0000000000000000;
        memory[266] = 16'b0000000000000000;
        memory[267] = 16'b0000000000000000;
        memory[268] = 16'b0000000000000000;
        memory[269] = 16'b0000000000000000;
        memory[270] = 16'b0000000000000000;
        memory[271] = 16'b0000000000000000;

        // Flat symbol (♭) starting at address 
        memory[272] = 16'b0000000000000000;
        memory[273] = 16'b0000000100000000;
        memory[274] = 16'b0000001100000000;
        memory[275] = 16'b0000001100000000;
        memory[276] = 16'b0000001100000000;
        memory[277] = 16'b0000001111111100;
        memory[278] = 16'b0000001100000110;
        memory[279] = 16'b0000001100000110;
        memory[280] = 16'b0000001100000110;
        memory[281] = 16'b0000001111111100;
        memory[282] = 16'b0000000000000000;
        memory[283] = 16'b0000000000000000;
        memory[284] = 16'b0000000000000000;
        memory[285] = 16'b0000000000000000;
        memory[286] = 16'b0000000000000000;
        memory[287] = 16'b0000000000000000;

    end

    always @(posedge clk_in ) begin
        data <= memory[addr]; // Output the 16-bit row at the given address
    end

endmodule