module NoteLoader(
    input logic clk_in,                     // Clock signal
    input logic rst_in,                   // rst_in signal
    input wire start,
    output logic [15:0] results [31:0],  // Array to store 32 results
    output logic done                    // Signal indicating processing is complete
);

    // Simulated BRAM (for testing or FPGA instantiation)
    logic [7:0] bram [0:64000];    // 512x16 BRAM storage

    // always_comb begin
//         bram[0] = 127;
// bram[1] = 140;
// bram[2] = 152;
// bram[3] = 165;
// bram[4] = 177;
// bram[5] = 189;
// bram[6] = 200;
// bram[7] = 210;
// bram[8] = 220;
// bram[9] = 228;
// bram[10] = 235;
// bram[11] = 241;
// bram[12] = 246;
// bram[13] = 250;
// bram[14] = 252;
// bram[15] = 253;
// bram[16] = 253;
// bram[17] = 251;
// bram[18] = 249;
// bram[19] = 244;
// bram[20] = 239;
// bram[21] = 232;
// bram[22] = 224;
// bram[23] = 215;
// bram[24] = 206;
// bram[25] = 195;
// bram[26] = 184;
// bram[27] = 172;
// bram[28] = 159;
// bram[29] = 146;
// bram[30] = 133;
// bram[31] = 120;
// bram[32] = 107;
// bram[33] = 95;
// bram[34] = 82;
// bram[35] = 70;
// bram[36] = 59;
// bram[37] = 48;
// bram[38] = 38;
// bram[39] = 29;
// bram[40] = 21;
// bram[41] = 15;
// bram[42] = 9;
// bram[43] = 5;
// bram[44] = 2;
// bram[45] = 0;
// bram[46] = 0;
// bram[47] = 0;
// bram[48] = 3;
// bram[49] = 6;
// bram[50] = 11;
// bram[51] = 17;
// bram[52] = 24;
// bram[53] = 33;
// bram[54] = 42;
// bram[55] = 52;
// bram[56] = 63;
// bram[57] = 75;
// bram[58] = 87;
// bram[59] = 100;
// bram[60] = 113;
// bram[61] = 126;
// bram[62] = 139;
// bram[63] = 152;
// bram[64] = 164;
// bram[65] = 176;
// bram[66] = 188;
// bram[67] = 199;
// bram[68] = 210;
// bram[69] = 219;
// bram[70] = 227;
// bram[71] = 235;
// bram[72] = 241;
// bram[73] = 246;
// bram[74] = 250;
// bram[75] = 252;
// bram[76] = 253;
// bram[77] = 253;
// bram[78] = 252;
// bram[79] = 249;
// bram[80] = 245;
// bram[81] = 239;
// bram[82] = 233;
// bram[83] = 225;
// bram[84] = 216;
// bram[85] = 206;
// bram[86] = 196;
// bram[87] = 184;
// bram[88] = 173;
// bram[89] = 160;
// bram[90] = 147;
// bram[91] = 134;
// bram[92] = 121;
// bram[93] = 108;
// bram[94] = 95;
// bram[95] = 83;
// bram[96] = 71;
// bram[97] = 60;
// bram[98] = 49;
// bram[99] = 39;
// bram[100] = 30;
// bram[101] = 22;
// bram[102] = 15;
// bram[103] = 9;
// bram[104] = 5;
// bram[105] = 2;
// bram[106] = 0;
// bram[107] = 0;
// bram[108] = 0;
// bram[109] = 3;
// bram[110] = 6;
// bram[111] = 11;
// bram[112] = 17;
// bram[113] = 24;
// bram[114] = 32;
// bram[115] = 41;
// bram[116] = 52;
// bram[117] = 62;
// bram[118] = 74;
// bram[119] = 86;
// bram[120] = 99;
// bram[121] = 112;
// bram[122] = 125;
// bram[123] = 138;
// bram[124] = 151;
// bram[125] = 163;
// bram[126] = 176;
// bram[127] = 187;
// bram[128] = 199;
// bram[129] = 209;
// bram[130] = 218;
// bram[131] = 227;
// bram[132] = 234;
// bram[133] = 241;
// bram[134] = 246;
// bram[135] = 250;
// bram[136] = 252;
// bram[137] = 253;
// bram[138] = 253;
// bram[139] = 252;
// bram[140] = 249;
// bram[141] = 245;
// bram[142] = 240;
// bram[143] = 233;
// bram[144] = 225;
// bram[145] = 217;
// bram[146] = 207;
// bram[147] = 196;
// bram[148] = 185;
// bram[149] = 173;
// bram[150] = 161;
// bram[151] = 148;
// bram[152] = 135;
// bram[153] = 122;
// bram[154] = 109;
// bram[155] = 96;
// bram[156] = 84;
// bram[157] = 72;
// bram[158] = 60;
// bram[159] = 50;
// bram[160] = 40;
// bram[161] = 31;
// bram[162] = 22;
// bram[163] = 16;
// bram[164] = 10;
// bram[165] = 5;
// bram[166] = 2;
// bram[167] = 0;
// bram[168] = 0;
// bram[169] = 0;
// bram[170] = 2;
// bram[171] = 6;
// bram[172] = 10;
// bram[173] = 16;
// bram[174] = 23;
// bram[175] = 32;
// bram[176] = 41;
// bram[177] = 51;
// bram[178] = 62;
// bram[179] = 73;
// bram[180] = 85;
// bram[181] = 98;
// bram[182] = 111;
// bram[183] = 124;
// bram[184] = 137;
// bram[185] = 150;
// bram[186] = 163;
// bram[187] = 175;
// bram[188] = 187;
// bram[189] = 198;
// bram[190] = 208;
// bram[191] = 218;
// bram[192] = 226;
// bram[193] = 234;
// bram[194] = 240;
// bram[195] = 245;
// bram[196] = 249;
// bram[197] = 252;
// bram[198] = 253;
// bram[199] = 253;
// bram[200] = 252;
// bram[201] = 249;
// bram[202] = 245;
// bram[203] = 240;
// bram[204] = 234;
// bram[205] = 226;
// bram[206] = 217;
// bram[207] = 208;
// bram[208] = 197;
// bram[209] = 186;
// bram[210] = 174;
// bram[211] = 162;
// bram[212] = 149;
// bram[213] = 136;
// bram[214] = 123;
// bram[215] = 110;
// bram[216] = 97;
// bram[217] = 85;
// bram[218] = 73;
// bram[219] = 61;
// bram[220] = 50;
// bram[221] = 40;
// bram[222] = 31;
// bram[223] = 23;
// bram[224] = 16;
// bram[225] = 10;
// bram[226] = 6;
// bram[227] = 2;
// bram[228] = 0;
// bram[229] = 0;
// bram[230] = 0;
// bram[231] = 2;
// bram[232] = 5;
// bram[233] = 10;
// bram[234] = 16;
// bram[235] = 23;
// bram[236] = 31;
// bram[237] = 40;
// bram[238] = 50;
// bram[239] = 61;
// bram[240] = 72;
// bram[241] = 85;
// bram[242] = 97;
// bram[243] = 110;
// bram[244] = 123;
// bram[245] = 136;
// bram[246] = 149;
// bram[247] = 162;
// bram[248] = 174;
// bram[249] = 186;
// bram[250] = 197;
// bram[251] = 208;
// bram[252] = 217;
// bram[253] = 226;
// bram[254] = 233;
// bram[255] = 240;
// bram[256] = 245;
// bram[257] = 249;
// bram[258] = 252;
// bram[259] = 253;
// bram[260] = 253;
// bram[261] = 252;
// bram[262] = 249;
// bram[263] = 246;
// bram[264] = 240;
// bram[265] = 234;
// bram[266] = 226;
// bram[267] = 218;
// bram[268] = 208;
// bram[269] = 198;
// bram[270] = 187;
// bram[271] = 175;
// bram[272] = 163;
// bram[273] = 150;
// bram[274] = 137;
// bram[275] = 124;
// bram[276] = 111;
// bram[277] = 98;
// bram[278] = 86;
// bram[279] = 73;
// bram[280] = 62;
// bram[281] = 51;
// bram[282] = 41;
// bram[283] = 32;
// bram[284] = 24;
// bram[285] = 16;
// bram[286] = 11;
// bram[287] = 6;
// bram[288] = 2;
// bram[289] = 0;
// bram[290] = 0;
// bram[291] = 0;
// bram[292] = 2;
// bram[293] = 5;
// bram[294] = 10;
// bram[295] = 15;
// bram[296] = 22;
// bram[297] = 30;
// bram[298] = 39;
// bram[299] = 49;
// bram[300] = 60;
// bram[301] = 72;
// bram[302] = 84;
// bram[303] = 96;
// bram[304] = 109;
// bram[305] = 122;
// bram[306] = 135;
// bram[307] = 148;
// bram[308] = 161;
// bram[309] = 173;
// bram[310] = 185;
// bram[311] = 196;
// bram[312] = 207;
// bram[313] = 217;
// bram[314] = 225;
// bram[315] = 233;
// bram[316] = 239;
// bram[317] = 245;
// bram[318] = 249;
// bram[319] = 252;
// bram[320] = 253;
// bram[321] = 253;
// bram[322] = 252;
// bram[323] = 250;
// bram[324] = 246;
// bram[325] = 241;
// bram[326] = 234;
// bram[327] = 227;
// bram[328] = 219;
// bram[329] = 209;
// bram[330] = 199;
// bram[331] = 188;
// bram[332] = 176;
// bram[333] = 164;
// bram[334] = 151;
// bram[335] = 138;
// bram[336] = 125;
// bram[337] = 112;
// bram[338] = 99;
// bram[339] = 86;
// bram[340] = 74;
// bram[341] = 63;
// bram[342] = 52;
// bram[343] = 42;
// bram[344] = 32;
// bram[345] = 24;
// bram[346] = 17;
// bram[347] = 11;
// bram[348] = 6;
// bram[349] = 3;
// bram[350] = 0;
// bram[351] = 0;
// bram[352] = 0;
// bram[353] = 2;
// bram[354] = 5;
// bram[355] = 9;
// bram[356] = 15;
// bram[357] = 22;
// bram[358] = 30;
// bram[359] = 39;
// bram[360] = 49;
// bram[361] = 59;
// bram[362] = 71;
// bram[363] = 83;
// bram[364] = 95;
// bram[365] = 108;
// bram[366] = 121;
// bram[367] = 134;
// bram[368] = 147;
// bram[369] = 160;
// bram[370] = 172;
// bram[371] = 184;
// bram[372] = 196;
// bram[373] = 206;
// bram[374] = 216;
// bram[375] = 225;
// bram[376] = 232;
// bram[377] = 239;
// bram[378] = 245;
// bram[379] = 249;
// bram[380] = 252;
// bram[381] = 253;
// bram[382] = 253;
// bram[383] = 252;
// bram[384] = 250;
// bram[385] = 246;
// bram[386] = 241;
// bram[387] = 235;
// bram[388] = 228;
// bram[389] = 219;
// bram[390] = 210;
// bram[391] = 199;
// bram[392] = 188;
// bram[393] = 177;
// bram[394] = 164;
// bram[395] = 152;
// bram[396] = 139;
// bram[397] = 126;
// bram[398] = 113;
// bram[399] = 100;
// bram[400] = 87;
// bram[401] = 75;
// bram[402] = 63;
// bram[403] = 52;
// bram[404] = 42;
// bram[405] = 33;
// bram[406] = 25;
// bram[407] = 17;
// bram[408] = 11;
// bram[409] = 6;
// bram[410] = 3;
// bram[411] = 0;
// bram[412] = 0;
// bram[413] = 0;
// bram[414] = 2;
// bram[415] = 5;
// bram[416] = 9;
// bram[417] = 15;
// bram[418] = 21;
// bram[419] = 29;
// bram[420] = 38;
// bram[421] = 48;
// bram[422] = 59;
// bram[423] = 70;
// bram[424] = 82;
// bram[425] = 94;
// bram[426] = 107;
// bram[427] = 120;
// bram[428] = 133;
// bram[429] = 146;
// bram[430] = 159;
// bram[431] = 171;
// bram[432] = 183;
// bram[433] = 195;
// bram[434] = 205;
// bram[435] = 215;
// bram[436] = 224;
// bram[437] = 232;
// bram[438] = 239;
// bram[439] = 244;
// bram[440] = 248;
// bram[441] = 251;
// bram[442] = 253;
// bram[443] = 253;
// bram[444] = 252;
// bram[445] = 250;
// bram[446] = 246;
// bram[447] = 242;
// bram[448] = 235;
// bram[449] = 228;
// bram[450] = 220;
// bram[451] = 210;
// bram[452] = 200;
// bram[453] = 189;
// bram[454] = 177;
// bram[455] = 165;
// bram[456] = 153;
// bram[457] = 140;
// bram[458] = 127;
// bram[459] = 114;
// bram[460] = 101;
// bram[461] = 88;
// bram[462] = 76;
// bram[463] = 64;
// bram[464] = 53;
// bram[465] = 43;
// bram[466] = 34;
// bram[467] = 25;
// bram[468] = 18;
// bram[469] = 12;
// bram[470] = 7;
// bram[471] = 3;
// bram[472] = 1;
// bram[473] = 0;
// bram[474] = 0;
// bram[475] = 1;
// bram[476] = 4;
// bram[477] = 9;
// bram[478] = 14;
// bram[479] = 21;
// bram[480] = 29;
// bram[481] = 37;
// bram[482] = 47;
// bram[483] = 58;
// bram[484] = 69;
// bram[485] = 81;
// bram[486] = 94;
// bram[487] = 106;
// bram[488] = 119;
// bram[489] = 132;
// bram[490] = 145;
// bram[491] = 158;
// bram[492] = 171;
// bram[493] = 183;
// bram[494] = 194;
// bram[495] = 205;
// bram[496] = 215;
// bram[497] = 224;
// bram[498] = 231;
// bram[499] = 238;
// bram[500] = 244;
// bram[501] = 248;
// bram[502] = 251;
// bram[503] = 253;
// bram[504] = 253;
// bram[505] = 253;
// bram[506] = 250;
// bram[507] = 247;
// bram[508] = 242;
// bram[509] = 236;
// bram[510] = 229;
// bram[511] = 220;
// bram[512] = 211;
// bram[513] = 201;
// bram[514] = 190;
// bram[515] = 178;
// bram[516] = 166;
// bram[517] = 154;
// bram[518] = 141;
// bram[519] = 128;
// bram[520] = 115;
// bram[521] = 102;
// bram[522] = 89;
// bram[523] = 77;
// bram[524] = 65;
// bram[525] = 54;
// bram[526] = 44;
// bram[527] = 34;
// bram[528] = 26;
// bram[529] = 18;
// bram[530] = 12;
// bram[531] = 7;
// bram[532] = 3;
// bram[533] = 1;
// bram[534] = 0;
// bram[535] = 0;
// bram[536] = 1;
// bram[537] = 4;
// bram[538] = 8;
// bram[539] = 14;
// bram[540] = 20;
// bram[541] = 28;
// bram[542] = 37;
// bram[543] = 47;
// bram[544] = 57;
// bram[545] = 68;
// bram[546] = 80;
// bram[547] = 93;
// bram[548] = 105;
// bram[549] = 118;
// bram[550] = 131;
// bram[551] = 144;
// bram[552] = 157;
// bram[553] = 170;
// bram[554] = 182;
// bram[555] = 193;
// bram[556] = 204;
// bram[557] = 214;
// bram[558] = 223;
// bram[559] = 231;
// bram[560] = 238;
// bram[561] = 243;
// bram[562] = 248;
// bram[563] = 251;
// bram[564] = 253;
// bram[565] = 253;
// bram[566] = 253;
// bram[567] = 251;
// bram[568] = 247;
// bram[569] = 242;
// bram[570] = 236;
// bram[571] = 229;
// bram[572] = 221;
// bram[573] = 212;
// bram[574] = 202;
// bram[575] = 191;
// bram[576] = 179;
// bram[577] = 167;
// bram[578] = 154;
// bram[579] = 142;
// bram[580] = 128;
// bram[581] = 115;
// bram[582] = 103;
// bram[583] = 90;
// bram[584] = 78;
// bram[585] = 66;
// bram[586] = 55;
// bram[587] = 44;
// bram[588] = 35;
// bram[589] = 26;
// bram[590] = 19;
// bram[591] = 12;
// bram[592] = 7;
// bram[593] = 3;
// bram[594] = 1;
// bram[595] = 0;
// bram[596] = 0;
// bram[597] = 1;
// bram[598] = 4;
// bram[599] = 8;
// bram[600] = 13;
// bram[601] = 20;
// bram[602] = 28;
// bram[603] = 36;
// bram[604] = 46;
// bram[605] = 56;
// bram[606] = 68;
// bram[607] = 79;
// bram[608] = 92;
// bram[609] = 105;
// bram[610] = 118;
// bram[611] = 131;
// bram[612] = 144;
// bram[613] = 156;
// bram[614] = 169;
// bram[615] = 181;
// bram[616] = 193;
// bram[617] = 203;
// bram[618] = 213;
// bram[619] = 222;
// bram[620] = 230;
// bram[621] = 237;
// bram[622] = 243;
// bram[623] = 248;
// bram[624] = 251;
// bram[625] = 253;
// bram[626] = 253;
// bram[627] = 253;
// bram[628] = 251;
// bram[629] = 247;
// bram[630] = 243;
// bram[631] = 237;
// bram[632] = 230;
// bram[633] = 222;
// bram[634] = 212;
// bram[635] = 202;
// bram[636] = 191;
// bram[637] = 180;
// bram[638] = 168;
// bram[639] = 155;
// bram[640] = 142;
// bram[641] = 129;
// bram[642] = 116;
// bram[643] = 103;
// bram[644] = 91;
// bram[645] = 78;
// bram[646] = 67;
// bram[647] = 55;
// bram[648] = 45;
// bram[649] = 35;
// bram[650] = 27;
// bram[651] = 19;
// bram[652] = 13;
// bram[653] = 8;
// bram[654] = 4;
// bram[655] = 1;
// bram[656] = 0;
// bram[657] = 0;
// bram[658] = 1;
// bram[659] = 4;
// bram[660] = 8;
// bram[661] = 13;
// bram[662] = 19;
// bram[663] = 27;
// bram[664] = 36;
// bram[665] = 45;
// bram[666] = 56;
// bram[667] = 67;
// bram[668] = 79;
// bram[669] = 91;
// bram[670] = 104;
// bram[671] = 117;
// bram[672] = 130;
// bram[673] = 143;
// bram[674] = 156;
// bram[675] = 168;
// bram[676] = 180;
// bram[677] = 192;
// bram[678] = 203;
// bram[679] = 213;
// bram[680] = 222;
// bram[681] = 230;
// bram[682] = 237;
// bram[683] = 243;
// bram[684] = 247;
// bram[685] = 251;
// bram[686] = 253;
// bram[687] = 253;
// bram[688] = 253;
// bram[689] = 251;
// bram[690] = 248;
// bram[691] = 243;
// bram[692] = 237;
// bram[693] = 230;
// bram[694] = 222;
// bram[695] = 213;
// bram[696] = 203;
// bram[697] = 192;
// bram[698] = 181;
// bram[699] = 169;
// bram[700] = 156;
// bram[701] = 143;
// bram[702] = 130;
// bram[703] = 117;
// bram[704] = 104;
// bram[705] = 92;
// bram[706] = 79;
// bram[707] = 67;
// bram[708] = 56;
// bram[709] = 46;
// bram[710] = 36;
// bram[711] = 27;
// bram[712] = 20;
// bram[713] = 13;
// bram[714] = 8;
// bram[715] = 4;
// bram[716] = 1;
// bram[717] = 0;
// bram[718] = 0;
// bram[719] = 1;
// bram[720] = 3;
// bram[721] = 7;
// bram[722] = 13;
// bram[723] = 19;
// bram[724] = 26;
// bram[725] = 35;
// bram[726] = 44;
// bram[727] = 55;
// bram[728] = 66;
// bram[729] = 78;
// bram[730] = 90;
// bram[731] = 103;
// bram[732] = 116;
// bram[733] = 129;
// bram[734] = 142;
// bram[735] = 155;
// bram[736] = 167;
// bram[737] = 179;
// bram[738] = 191;
// bram[739] = 202;
// bram[740] = 212;
// bram[741] = 221;
// bram[742] = 229;
// bram[743] = 236;
// bram[744] = 242;
// bram[745] = 247;
// bram[746] = 251;
// bram[747] = 253;
// bram[748] = 253;
// bram[749] = 253;
// bram[750] = 251;
// bram[751] = 248;
// bram[752] = 243;
// bram[753] = 238;
// bram[754] = 231;
// bram[755] = 223;
// bram[756] = 214;
// bram[757] = 204;
// bram[758] = 193;
// bram[759] = 182;
// bram[760] = 170;
// bram[761] = 157;
// bram[762] = 144;
// bram[763] = 131;
// bram[764] = 118;
// bram[765] = 105;
// bram[766] = 92;
// bram[767] = 80;
// bram[768] = 68;
// bram[769] = 57;
// bram[770] = 46;
// bram[771] = 37;
// bram[772] = 28;
// bram[773] = 20;
// bram[774] = 14;
// bram[775] = 8;
// bram[776] = 4;
// bram[777] = 1;
// bram[778] = 0;
// bram[779] = 0;
// bram[780] = 1;
// bram[781] = 3;
// bram[782] = 7;
// bram[783] = 12;
// bram[784] = 18;
// bram[785] = 26;
// bram[786] = 34;
// bram[787] = 44;
// bram[788] = 54;
// bram[789] = 65;
// bram[790] = 77;
// bram[791] = 89;
// bram[792] = 102;
// bram[793] = 115;
// bram[794] = 128;
// bram[795] = 141;
// bram[796] = 154;
// bram[797] = 166;
// bram[798] = 179;
// bram[799] = 190;
// bram[800] = 201;
// bram[801] = 211;
// bram[802] = 221;
// bram[803] = 229;
// bram[804] = 236;
// bram[805] = 242;
// bram[806] = 247;
// bram[807] = 250;
// bram[808] = 253;
// bram[809] = 253;
// bram[810] = 253;
// bram[811] = 251;
// bram[812] = 248;
// bram[813] = 244;
// bram[814] = 238;
// bram[815] = 231;
// bram[816] = 223;
// bram[817] = 214;
// bram[818] = 204;
// bram[819] = 194;
// bram[820] = 182;
// bram[821] = 170;
// bram[822] = 158;
// bram[823] = 145;
// bram[824] = 132;
// bram[825] = 119;
// bram[826] = 106;
// bram[827] = 93;
// bram[828] = 81;
// bram[829] = 69;
// bram[830] = 58;
// bram[831] = 47;
// bram[832] = 37;
// bram[833] = 28;
// bram[834] = 21;
// bram[835] = 14;
// bram[836] = 9;
// bram[837] = 4;
// bram[838] = 1;
// bram[839] = 0;
// bram[840] = 0;
// bram[841] = 1;
// bram[842] = 3;
// bram[843] = 7;
// bram[844] = 12;
// bram[845] = 18;
// bram[846] = 25;
// bram[847] = 34;
// bram[848] = 43;
// bram[849] = 53;
// bram[850] = 64;
// bram[851] = 76;
// bram[852] = 88;
// bram[853] = 101;
// bram[854] = 114;
// bram[855] = 127;
// bram[856] = 140;
// bram[857] = 153;
// bram[858] = 166;
// bram[859] = 178;
// bram[860] = 189;
// bram[861] = 200;
// bram[862] = 211;
// bram[863] = 220;
// bram[864] = 228;
// bram[865] = 236;
// bram[866] = 242;
// bram[867] = 247;
// bram[868] = 250;
// bram[869] = 252;
// bram[870] = 253;
// bram[871] = 253;
// bram[872] = 251;
// bram[873] = 248;
// bram[874] = 244;
// bram[875] = 239;
// bram[876] = 232;
// bram[877] = 224;
// bram[878] = 215;
// bram[879] = 205;
// bram[880] = 195;
// bram[881] = 183;
// bram[882] = 171;
// bram[883] = 159;
// bram[884] = 146;
// bram[885] = 133;
// bram[886] = 120;
// bram[887] = 107;
// bram[888] = 94;
// bram[889] = 82;
// bram[890] = 70;
// bram[891] = 58;
// bram[892] = 48;
// bram[893] = 38;
// bram[894] = 29;
// bram[895] = 21;
// bram[896] = 14;
// bram[897] = 9;
// bram[898] = 5;
// bram[899] = 2;
// bram[900] = 0;
// bram[901] = 0;
// bram[902] = 1;
// bram[903] = 3;
// bram[904] = 6;
// bram[905] = 11;
// bram[906] = 17;
// bram[907] = 25;
// bram[908] = 33;
// bram[909] = 42;
// bram[910] = 53;
// bram[911] = 64;
// bram[912] = 75;
// bram[913] = 88;
// bram[914] = 100;
// bram[915] = 113;
// bram[916] = 126;
// bram[917] = 139;
// bram[918] = 152;
// bram[919] = 165;
// bram[920] = 177;
// bram[921] = 189;
// bram[922] = 200;
// bram[923] = 210;
// bram[924] = 219;
// bram[925] = 228;
// bram[926] = 235;
// bram[927] = 241;
// bram[928] = 246;
// bram[929] = 250;
// bram[930] = 252;
// bram[931] = 253;
// bram[932] = 253;
// bram[933] = 252;
// bram[934] = 249;
// bram[935] = 244;
// bram[936] = 239;
// bram[937] = 232;
// bram[938] = 224;
// bram[939] = 216;
// bram[940] = 206;
// bram[941] = 195;
// bram[942] = 184;
// bram[943] = 172;
// bram[944] = 160;
// bram[945] = 147;
// bram[946] = 134;
// bram[947] = 121;
// bram[948] = 108;
// bram[949] = 95;
// bram[950] = 83;
// bram[951] = 71;
// bram[952] = 59;
// bram[953] = 48;
// bram[954] = 39;
// bram[955] = 30;
// bram[956] = 22;
// bram[957] = 15;
// bram[958] = 9;
// bram[959] = 5;
// bram[960] = 2;
// bram[961] = 0;
// bram[962] = 0;
// bram[963] = 0;
// bram[964] = 3;
// bram[965] = 6;
// bram[966] = 11;
// bram[967] = 17;
// bram[968] = 24;
// bram[969] = 32;
// bram[970] = 42;
// bram[971] = 52;
// bram[972] = 63;
// bram[973] = 75;
// bram[974] = 87;
// bram[975] = 99;
// bram[976] = 112;
// bram[977] = 125;
// bram[978] = 138;
// bram[979] = 151;
// bram[980] = 164;
// bram[981] = 176;
// bram[982] = 188;
// bram[983] = 199;
// bram[984] = 209;
// bram[985] = 219;
// bram[986] = 227;
// bram[987] = 235;
// bram[988] = 241;
// bram[989] = 246;
// bram[990] = 250;
// bram[991] = 252;
// bram[992] = 253;
// bram[993] = 253;
// bram[994] = 252;
// bram[995] = 249;
// bram[996] = 245;
// bram[997] = 239;
// bram[998] = 233;
// bram[999] = 225;
// bram[1000] = 216;
// bram[1001] = 207;
// bram[1002] = 196;
// bram[1003] = 185;
// bram[1004] = 173;
// bram[1005] = 160;
// bram[1006] = 148;
// bram[1007] = 135;
// bram[1008] = 122;
// bram[1009] = 109;
// bram[1010] = 96;
// bram[1011] = 83;
// bram[1012] = 71;
// bram[1013] = 60;
// bram[1014] = 49;
// bram[1015] = 39;
// bram[1016] = 30;
// bram[1017] = 22;
// bram[1018] = 15;
// bram[1019] = 10;
// bram[1020] = 5;
// bram[1021] = 2;
// bram[1022] = 0;
// bram[1023] = 0;
// bram[1024] = 0;
// bram[1025] = 2;
// bram[1026] = 6;
// bram[1027] = 11;
// bram[1028] = 17;
// bram[1029] = 24;
// bram[1030] = 32;
// bram[1031] = 41;
// bram[1032] = 51;
// bram[1033] = 62;
// bram[1034] = 74;
// bram[1035] = 86;
// bram[1036] = 98;
// bram[1037] = 111;
// bram[1038] = 124;
// bram[1039] = 137;
// bram[1040] = 150;
// bram[1041] = 163;
// bram[1042] = 175;
// bram[1043] = 187;
// bram[1044] = 198;
// bram[1045] = 209;
// bram[1046] = 218;
// bram[1047] = 227;
// bram[1048] = 234;
// bram[1049] = 241;
// bram[1050] = 246;
// bram[1051] = 250;
// bram[1052] = 252;
// bram[1053] = 253;
// bram[1054] = 253;
// bram[1055] = 252;
// bram[1056] = 249;
// bram[1057] = 245;
// bram[1058] = 240;
// bram[1059] = 233;
// bram[1060] = 226;
// bram[1061] = 217;
// bram[1062] = 207;
// bram[1063] = 197;
// bram[1064] = 186;
// bram[1065] = 174;
// bram[1066] = 161;
// bram[1067] = 149;
// bram[1068] = 136;
// bram[1069] = 123;
// bram[1070] = 110;
// bram[1071] = 97;
// bram[1072] = 84;
// bram[1073] = 72;
// bram[1074] = 61;
// bram[1075] = 50;
// bram[1076] = 40;
// bram[1077] = 31;
// bram[1078] = 23;
// bram[1079] = 16;
// bram[1080] = 10;
// bram[1081] = 5;
// bram[1082] = 2;
// bram[1083] = 0;
// bram[1084] = 0;
// bram[1085] = 0;
// bram[1086] = 2;
// bram[1087] = 6;
// bram[1088] = 10;
// bram[1089] = 16;
// bram[1090] = 23;
// bram[1091] = 31;
// bram[1092] = 40;
// bram[1093] = 50;
// bram[1094] = 61;
// bram[1095] = 73;
// bram[1096] = 85;
// bram[1097] = 98;
// bram[1098] = 110;
// bram[1099] = 123;
// bram[1100] = 136;
// bram[1101] = 149;
// bram[1102] = 162;
// bram[1103] = 174;
// bram[1104] = 186;
// bram[1105] = 197;
// bram[1106] = 208;
// bram[1107] = 217;
// bram[1108] = 226;
// bram[1109] = 234;
// bram[1110] = 240;
// bram[1111] = 245;
// bram[1112] = 249;
// bram[1113] = 252;
// bram[1114] = 253;
// bram[1115] = 253;
// bram[1116] = 252;
// bram[1117] = 249;
// bram[1118] = 245;
// bram[1119] = 240;
// bram[1120] = 234;
// bram[1121] = 226;
// bram[1122] = 218;
// bram[1123] = 208;
// bram[1124] = 198;
// bram[1125] = 186;
// bram[1126] = 175;
// bram[1127] = 162;
// bram[1128] = 150;
// bram[1129] = 137;
// bram[1130] = 124;
// bram[1131] = 110;
// bram[1132] = 98;
// bram[1133] = 85;
// bram[1134] = 73;
// bram[1135] = 61;
// bram[1136] = 51;
// bram[1137] = 41;
// bram[1138] = 31;
// bram[1139] = 23;
// bram[1140] = 16;
// bram[1141] = 10;
// bram[1142] = 6;
// bram[1143] = 2;
// bram[1144] = 0;
// bram[1145] = 0;
// bram[1146] = 0;
// bram[1147] = 2;
// bram[1148] = 5;
// bram[1149] = 10;
// bram[1150] = 16;
// bram[1151] = 23;
// bram[1152] = 31;
// bram[1153] = 40;
// bram[1154] = 50;
// bram[1155] = 61;
// bram[1156] = 72;
// bram[1157] = 84;
// bram[1158] = 97;
// bram[1159] = 109;
// bram[1160] = 123;
// bram[1161] = 136;
// bram[1162] = 149;
// bram[1163] = 161;
// bram[1164] = 174;
// bram[1165] = 185;
// bram[1166] = 197;
// bram[1167] = 207;
// bram[1168] = 217;
// bram[1169] = 226;
// bram[1170] = 233;
// bram[1171] = 240;
// bram[1172] = 245;
// bram[1173] = 249;
// bram[1174] = 252;
// bram[1175] = 253;
// bram[1176] = 253;
// bram[1177] = 252;
// bram[1178] = 250;
// bram[1179] = 246;
// bram[1180] = 241;
// bram[1181] = 234;
// bram[1182] = 227;
// bram[1183] = 218;
// bram[1184] = 209;
// bram[1185] = 198;
// bram[1186] = 187;
// bram[1187] = 175;
// bram[1188] = 163;
// bram[1189] = 150;
// bram[1190] = 137;
// bram[1191] = 124;
// bram[1192] = 111;
// bram[1193] = 99;
// bram[1194] = 86;
// bram[1195] = 74;
// bram[1196] = 62;
// bram[1197] = 51;
// bram[1198] = 41;
// bram[1199] = 32;
// bram[1200] = 24;
// bram[1201] = 17;
// bram[1202] = 11;
// bram[1203] = 6;
// bram[1204] = 2;
// bram[1205] = 0;
// bram[1206] = 0;
// bram[1207] = 0;
// bram[1208] = 2;
// bram[1209] = 5;
// bram[1210] = 10;
// bram[1211] = 15;
// bram[1212] = 22;
// bram[1213] = 30;
// bram[1214] = 39;
// bram[1215] = 49;
// bram[1216] = 60;
// bram[1217] = 71;
// bram[1218] = 83;
// bram[1219] = 96;
// bram[1220] = 109;
// bram[1221] = 122;
// bram[1222] = 135;
// bram[1223] = 148;
// bram[1224] = 160;
// bram[1225] = 173;
// bram[1226] = 185;
// bram[1227] = 196;
// bram[1228] = 207;
// bram[1229] = 216;
// bram[1230] = 225;
// bram[1231] = 233;
// bram[1232] = 239;
// bram[1233] = 245;
// bram[1234] = 249;
// bram[1235] = 252;
// bram[1236] = 253;
// bram[1237] = 253;
// bram[1238] = 252;
// bram[1239] = 250;
// bram[1240] = 246;
// bram[1241] = 241;
// bram[1242] = 235;
// bram[1243] = 227;
// bram[1244] = 219;
// bram[1245] = 209;
// bram[1246] = 199;
// bram[1247] = 188;
// bram[1248] = 176;
// bram[1249] = 164;
// bram[1250] = 151;
// bram[1251] = 138;
// bram[1252] = 125;
// bram[1253] = 112;
// bram[1254] = 99;
// bram[1255] = 87;
// bram[1256] = 75;
// bram[1257] = 63;
// bram[1258] = 52;
// bram[1259] = 42;
// bram[1260] = 33;
// bram[1261] = 24;
// bram[1262] = 17;
// bram[1263] = 11;
// bram[1264] = 6;
// bram[1265] = 3;
// bram[1266] = 0;
// bram[1267] = 0;
// bram[1268] = 0;
// bram[1269] = 2;
// bram[1270] = 5;
// bram[1271] = 9;
// bram[1272] = 15;
// bram[1273] = 22;
// bram[1274] = 30;
// bram[1275] = 38;
// bram[1276] = 48;
// bram[1277] = 59;
// bram[1278] = 70;
// bram[1279] = 82;
// bram[1280] = 95;
// bram[1281] = 108;
// bram[1282] = 121;
// bram[1283] = 134;
// bram[1284] = 147;
// bram[1285] = 160;
// bram[1286] = 172;
// bram[1287] = 184;
// bram[1288] = 195;
// bram[1289] = 206;
// bram[1290] = 216;
// bram[1291] = 224;
// bram[1292] = 232;
// bram[1293] = 239;
// bram[1294] = 244;
// bram[1295] = 249;
// bram[1296] = 252;
// bram[1297] = 253;
// bram[1298] = 253;
// bram[1299] = 252;
// bram[1300] = 250;
// bram[1301] = 246;
// bram[1302] = 241;
// bram[1303] = 235;
// bram[1304] = 228;
// bram[1305] = 219;
// bram[1306] = 210;
// bram[1307] = 200;
// bram[1308] = 189;
// bram[1309] = 177;
// bram[1310] = 165;
// bram[1311] = 152;
// bram[1312] = 139;
// bram[1313] = 126;
// bram[1314] = 113;
// bram[1315] = 100;
// bram[1316] = 88;
// bram[1317] = 75;
// bram[1318] = 64;
// bram[1319] = 53;
// bram[1320] = 43;
// bram[1321] = 33;
// bram[1322] = 25;
// bram[1323] = 18;
// bram[1324] = 11;
// bram[1325] = 7;
// bram[1326] = 3;
// bram[1327] = 1;
// bram[1328] = 0;
// bram[1329] = 0;
// bram[1330] = 2;
// bram[1331] = 5;
// bram[1332] = 9;
// bram[1333] = 14;
// bram[1334] = 21;
// bram[1335] = 29;
// bram[1336] = 38;
// bram[1337] = 48;
// bram[1338] = 58;
// bram[1339] = 70;
// bram[1340] = 82;
// bram[1341] = 94;
// bram[1342] = 107;
// bram[1343] = 120;
// bram[1344] = 133;
// bram[1345] = 146;
// bram[1346] = 159;
// bram[1347] = 171;
// bram[1348] = 183;
// bram[1349] = 194;
// bram[1350] = 205;
// bram[1351] = 215;
// bram[1352] = 224;
// bram[1353] = 232;
// bram[1354] = 238;
// bram[1355] = 244;
// bram[1356] = 248;
// bram[1357] = 251;
// bram[1358] = 253;
// bram[1359] = 253;
// bram[1360] = 252;
// bram[1361] = 250;
// bram[1362] = 247;
// bram[1363] = 242;
// bram[1364] = 236;
// bram[1365] = 228;
// bram[1366] = 220;
// bram[1367] = 211;
// bram[1368] = 201;
// bram[1369] = 190;
// bram[1370] = 178;
// bram[1371] = 166;
// bram[1372] = 153;
// bram[1373] = 140;
// bram[1374] = 127;
// bram[1375] = 114;
// bram[1376] = 101;
// bram[1377] = 88;
// bram[1378] = 76;
// bram[1379] = 65;
// bram[1380] = 53;
// bram[1381] = 43;
// bram[1382] = 34;
// bram[1383] = 25;
// bram[1384] = 18;
// bram[1385] = 12;
// bram[1386] = 7;
// bram[1387] = 3;
// bram[1388] = 1;
// bram[1389] = 0;
// bram[1390] = 0;
// bram[1391] = 1;
// bram[1392] = 4;
// bram[1393] = 9;
// bram[1394] = 14;
// bram[1395] = 21;
// bram[1396] = 28;
// bram[1397] = 37;
// bram[1398] = 47;
// bram[1399] = 58;
// bram[1400] = 69;
// bram[1401] = 81;
// bram[1402] = 93;
// bram[1403] = 106;
// bram[1404] = 119;
// bram[1405] = 132;
// bram[1406] = 145;
// bram[1407] = 158;
// bram[1408] = 170;
// bram[1409] = 182;
// bram[1410] = 194;
// bram[1411] = 204;
// bram[1412] = 214;
// bram[1413] = 223;
// bram[1414] = 231;
// bram[1415] = 238;
// bram[1416] = 244;
// bram[1417] = 248;
// bram[1418] = 251;
// bram[1419] = 253;
// bram[1420] = 253;
// bram[1421] = 253;
// bram[1422] = 250;
// bram[1423] = 247;
// bram[1424] = 242;
// bram[1425] = 236;
// bram[1426] = 229;
// bram[1427] = 221;
// bram[1428] = 211;
// bram[1429] = 201;
// bram[1430] = 190;
// bram[1431] = 179;
// bram[1432] = 167;
// bram[1433] = 154;
// bram[1434] = 141;
// bram[1435] = 128;
// bram[1436] = 115;
// bram[1437] = 102;
// bram[1438] = 89;
// bram[1439] = 77;
// bram[1440] = 65;
// bram[1441] = 54;
// bram[1442] = 44;
// bram[1443] = 34;
// bram[1444] = 26;
// bram[1445] = 18;
// bram[1446] = 12;
// bram[1447] = 7;
// bram[1448] = 3;
// bram[1449] = 1;
// bram[1450] = 0;
// bram[1451] = 0;
// bram[1452] = 1;
// bram[1453] = 4;
// bram[1454] = 8;
// bram[1455] = 14;
// bram[1456] = 20;
// bram[1457] = 28;
// bram[1458] = 37;
// bram[1459] = 46;
// bram[1460] = 57;
// bram[1461] = 68;
// bram[1462] = 80;
// bram[1463] = 92;
// bram[1464] = 105;
// bram[1465] = 118;
// bram[1466] = 131;
// bram[1467] = 144;
// bram[1468] = 157;
// bram[1469] = 169;
// bram[1470] = 181;
// bram[1471] = 193;
// bram[1472] = 204;
// bram[1473] = 214;
// bram[1474] = 223;
// bram[1475] = 231;
// bram[1476] = 238;
// bram[1477] = 243;
// bram[1478] = 248;
// bram[1479] = 251;
// bram[1480] = 253;
// bram[1481] = 253;
// bram[1482] = 253;
// bram[1483] = 251;
// bram[1484] = 247;
// bram[1485] = 242;
// bram[1486] = 237;
// bram[1487] = 229;
// bram[1488] = 221;
// bram[1489] = 212;
// bram[1490] = 202;
// bram[1491] = 191;
// bram[1492] = 179;
// bram[1493] = 167;
// bram[1494] = 155;
// bram[1495] = 142;
// bram[1496] = 129;
// bram[1497] = 116;
// bram[1498] = 103;
// bram[1499] = 90;
// bram[1500] = 78;
// bram[1501] = 66;
// bram[1502] = 55;
// bram[1503] = 45;
// bram[1504] = 35;
// bram[1505] = 26;
// bram[1506] = 19;
// bram[1507] = 13;
// bram[1508] = 7;
// bram[1509] = 4;
// bram[1510] = 1;
// bram[1511] = 0;
// bram[1512] = 0;
// bram[1513] = 1;
// bram[1514] = 4;
// bram[1515] = 8;
// bram[1516] = 13;
// bram[1517] = 20;
// bram[1518] = 27;
// bram[1519] = 36;
// bram[1520] = 46;
// bram[1521] = 56;
// bram[1522] = 67;
// bram[1523] = 79;
// bram[1524] = 91;
// bram[1525] = 104;
// bram[1526] = 117;
// bram[1527] = 130;
// bram[1528] = 143;
// bram[1529] = 156;
// bram[1530] = 169;
// bram[1531] = 181;
// bram[1532] = 192;
// bram[1533] = 203;
// bram[1534] = 213;
// bram[1535] = 222;
// bram[1536] = 230;
// bram[1537] = 237;
// bram[1538] = 243;
// bram[1539] = 248;
// bram[1540] = 251;
// bram[1541] = 253;
// bram[1542] = 253;
// bram[1543] = 253;
// bram[1544] = 251;
// bram[1545] = 247;
// bram[1546] = 243;
// bram[1547] = 237;
// bram[1548] = 230;
// bram[1549] = 222;
// bram[1550] = 213;
// bram[1551] = 203;
// bram[1552] = 192;
// bram[1553] = 180;
// bram[1554] = 168;
// bram[1555] = 156;
// bram[1556] = 143;
// bram[1557] = 130;
// bram[1558] = 117;
// bram[1559] = 104;
// bram[1560] = 91;
// bram[1561] = 79;
// bram[1562] = 67;
// bram[1563] = 56;
// bram[1564] = 45;
// bram[1565] = 36;
// bram[1566] = 27;
// bram[1567] = 19;
// bram[1568] = 13;
// bram[1569] = 8;
// bram[1570] = 4;
// bram[1571] = 1;
// bram[1572] = 0;
// bram[1573] = 0;
// bram[1574] = 1;
// bram[1575] = 4;
// bram[1576] = 8;
// bram[1577] = 13;
// bram[1578] = 19;
// bram[1579] = 27;
// bram[1580] = 35;
// bram[1581] = 45;
// bram[1582] = 55;
// bram[1583] = 66;
// bram[1584] = 78;
// bram[1585] = 91;
// bram[1586] = 103;
// bram[1587] = 116;
// bram[1588] = 129;
// bram[1589] = 142;
// bram[1590] = 155;
// bram[1591] = 168;
// bram[1592] = 180;
// bram[1593] = 191;
// bram[1594] = 202;
// bram[1595] = 212;
// bram[1596] = 221;
// bram[1597] = 230;
// bram[1598] = 237;
// bram[1599] = 243;
// bram[1600] = 247;
// bram[1601] = 251;
// bram[1602] = 253;
// bram[1603] = 253;
// bram[1604] = 253;
// bram[1605] = 251;
// bram[1606] = 248;
// bram[1607] = 243;
// bram[1608] = 237;
// bram[1609] = 230;
// bram[1610] = 222;
// bram[1611] = 213;
// bram[1612] = 203;
// bram[1613] = 193;
// bram[1614] = 181;
// bram[1615] = 169;
// bram[1616] = 157;
// bram[1617] = 144;
// bram[1618] = 131;
// bram[1619] = 118;
// bram[1620] = 105;
// bram[1621] = 92;
// bram[1622] = 80;
// bram[1623] = 68;
// bram[1624] = 56;
// bram[1625] = 46;
// bram[1626] = 36;
// bram[1627] = 28;
// bram[1628] = 20;
// bram[1629] = 13;
// bram[1630] = 8;
// bram[1631] = 4;
// bram[1632] = 1;
// bram[1633] = 0;
// bram[1634] = 0;
// bram[1635] = 1;
// bram[1636] = 3;
// bram[1637] = 7;
// bram[1638] = 12;
// bram[1639] = 19;
// bram[1640] = 26;
// bram[1641] = 35;
// bram[1642] = 44;
// bram[1643] = 55;
// bram[1644] = 66;
// bram[1645] = 77;
// bram[1646] = 90;
// bram[1647] = 102;
// bram[1648] = 115;
// bram[1649] = 128;
// bram[1650] = 141;
// bram[1651] = 154;
// bram[1652] = 167;
// bram[1653] = 179;
// bram[1654] = 191;
// bram[1655] = 202;
// bram[1656] = 212;
// bram[1657] = 221;
// bram[1658] = 229;
// bram[1659] = 236;
// bram[1660] = 242;
// bram[1661] = 247;
// bram[1662] = 250;
// bram[1663] = 253;
// bram[1664] = 253;
// bram[1665] = 253;
// bram[1666] = 251;
// bram[1667] = 248;
// bram[1668] = 244;
// bram[1669] = 238;
// bram[1670] = 231;
// bram[1671] = 223;
// bram[1672] = 214;
// bram[1673] = 204;
// bram[1674] = 193;
// bram[1675] = 182;
// bram[1676] = 170;
// bram[1677] = 157;
// bram[1678] = 145;
// bram[1679] = 132;
// bram[1680] = 119;
// bram[1681] = 106;
// bram[1682] = 93;
// bram[1683] = 80;
// bram[1684] = 68;
// bram[1685] = 57;
// bram[1686] = 47;
// bram[1687] = 37;
// bram[1688] = 28;
// bram[1689] = 20;
// bram[1690] = 14;
// bram[1691] = 8;
// bram[1692] = 4;
// bram[1693] = 1;
// bram[1694] = 0;
// bram[1695] = 0;
// bram[1696] = 1;
// bram[1697] = 3;
// bram[1698] = 7;
// bram[1699] = 12;
// bram[1700] = 18;
// bram[1701] = 26;
// bram[1702] = 34;
// bram[1703] = 43;
// bram[1704] = 54;
// bram[1705] = 65;
// bram[1706] = 77;
// bram[1707] = 89;
// bram[1708] = 102;
// bram[1709] = 114;
// bram[1710] = 127;
// bram[1711] = 141;
// bram[1712] = 153;
// bram[1713] = 166;
// bram[1714] = 178;
// bram[1715] = 190;
// bram[1716] = 201;
// bram[1717] = 211;
// bram[1718] = 220;
// bram[1719] = 229;
// bram[1720] = 236;
// bram[1721] = 242;
// bram[1722] = 247;
// bram[1723] = 250;
// bram[1724] = 253;
// bram[1725] = 253;
// bram[1726] = 253;
// bram[1727] = 251;
// bram[1728] = 248;
// bram[1729] = 244;
// bram[1730] = 238;
// bram[1731] = 231;
// bram[1732] = 224;
// bram[1733] = 215;
// bram[1734] = 205;
// bram[1735] = 194;
// bram[1736] = 183;
// bram[1737] = 171;
// bram[1738] = 158;
// bram[1739] = 145;
// bram[1740] = 132;
// bram[1741] = 119;
// bram[1742] = 106;
// bram[1743] = 94;
// bram[1744] = 81;
// bram[1745] = 69;
// bram[1746] = 58;
// bram[1747] = 47;
// bram[1748] = 38;
// bram[1749] = 29;
// bram[1750] = 21;
// bram[1751] = 14;
// bram[1752] = 9;
// bram[1753] = 4;
// bram[1754] = 1;
// bram[1755] = 0;
// bram[1756] = 0;
// bram[1757] = 1;
// bram[1758] = 3;
// bram[1759] = 7;
// bram[1760] = 12;
// bram[1761] = 18;
// bram[1762] = 25;
// bram[1763] = 33;
// bram[1764] = 43;
// bram[1765] = 53;
// bram[1766] = 64;
// bram[1767] = 76;
// bram[1768] = 88;
// bram[1769] = 101;
// bram[1770] = 114;
// bram[1771] = 127;
// bram[1772] = 140;
// bram[1773] = 153;
// bram[1774] = 165;
// bram[1775] = 177;
// bram[1776] = 189;
// bram[1777] = 200;
// bram[1778] = 210;
// bram[1779] = 220;
// bram[1780] = 228;
// bram[1781] = 235;
// bram[1782] = 241;
// bram[1783] = 246;
// bram[1784] = 250;
// bram[1785] = 252;
// bram[1786] = 253;
// bram[1787] = 253;
// bram[1788] = 251;
// bram[1789] = 248;
// bram[1790] = 244;
// bram[1791] = 239;
// bram[1792] = 232;
// bram[1793] = 224;
// bram[1794] = 215;
// bram[1795] = 206;
// bram[1796] = 195;
// bram[1797] = 184;
// bram[1798] = 172;
// bram[1799] = 159;
// bram[1800] = 146;
// bram[1801] = 133;
// bram[1802] = 120;
// bram[1803] = 107;
// bram[1804] = 95;
// bram[1805] = 82;
// bram[1806] = 70;
// bram[1807] = 59;
// bram[1808] = 48;
// bram[1809] = 38;
// bram[1810] = 29;
// bram[1811] = 21;
// bram[1812] = 15;
// bram[1813] = 9;
// bram[1814] = 5;
// bram[1815] = 2;
// bram[1816] = 0;
// bram[1817] = 0;
// bram[1818] = 0;
// bram[1819] = 3;
// bram[1820] = 6;
// bram[1821] = 11;
// bram[1822] = 17;
// bram[1823] = 25;
// bram[1824] = 33;
// bram[1825] = 42;
// bram[1826] = 52;
// bram[1827] = 63;
// bram[1828] = 75;
// bram[1829] = 87;
// bram[1830] = 100;
// bram[1831] = 113;
// bram[1832] = 126;
// bram[1833] = 139;
// bram[1834] = 152;
// bram[1835] = 164;
// bram[1836] = 177;
// bram[1837] = 188;
// bram[1838] = 199;
// bram[1839] = 210;
// bram[1840] = 219;
// bram[1841] = 228;
// bram[1842] = 235;
// bram[1843] = 241;
// bram[1844] = 246;
// bram[1845] = 250;
// bram[1846] = 252;
// bram[1847] = 253;
// bram[1848] = 253;
// bram[1849] = 252;
// bram[1850] = 249;
// bram[1851] = 245;
// bram[1852] = 239;
// bram[1853] = 232;
// bram[1854] = 225;
// bram[1855] = 216;
// bram[1856] = 206;
// bram[1857] = 196;
// bram[1858] = 184;
// bram[1859] = 172;
// bram[1860] = 160;
// bram[1861] = 147;
// bram[1862] = 134;
// bram[1863] = 121;
// bram[1864] = 108;
// bram[1865] = 95;
// bram[1866] = 83;
// bram[1867] = 71;
// bram[1868] = 59;
// bram[1869] = 49;
// bram[1870] = 39;
// bram[1871] = 30;
// bram[1872] = 22;
// bram[1873] = 15;
// bram[1874] = 9;
// bram[1875] = 5;
// bram[1876] = 2;
// bram[1877] = 0;
// bram[1878] = 0;
// bram[1879] = 0;
// bram[1880] = 3;
// bram[1881] = 6;
// bram[1882] = 11;
// bram[1883] = 17;
// bram[1884] = 24;
// bram[1885] = 32;
// bram[1886] = 41;
// bram[1887] = 52;
// bram[1888] = 63;
// bram[1889] = 74;
// bram[1890] = 86;
// bram[1891] = 99;
// bram[1892] = 112;
// bram[1893] = 125;
// bram[1894] = 138;
// bram[1895] = 151;
// bram[1896] = 163;
// bram[1897] = 176;
// bram[1898] = 188;
// bram[1899] = 199;
// bram[1900] = 209;
// bram[1901] = 218;
// bram[1902] = 227;
// bram[1903] = 234;
// bram[1904] = 241;
// bram[1905] = 246;
// bram[1906] = 250;
// bram[1907] = 252;
// bram[1908] = 253;
// bram[1909] = 253;
// bram[1910] = 252;
// bram[1911] = 249;
// bram[1912] = 245;
// bram[1913] = 240;
// bram[1914] = 233;
// bram[1915] = 225;
// bram[1916] = 217;
// bram[1917] = 207;
// bram[1918] = 196;
// bram[1919] = 185;
// bram[1920] = 173;
// bram[1921] = 161;
// bram[1922] = 148;
// bram[1923] = 135;
// bram[1924] = 122;
// bram[1925] = 109;
// bram[1926] = 96;
// bram[1927] = 84;
// bram[1928] = 72;
// bram[1929] = 60;
// bram[1930] = 49;
// bram[1931] = 39;
// bram[1932] = 30;
// bram[1933] = 22;
// bram[1934] = 15;
// bram[1935] = 10;
// bram[1936] = 5;
// bram[1937] = 2;
// bram[1938] = 0;
// bram[1939] = 0;
// bram[1940] = 0;
// bram[1941] = 2;
// bram[1942] = 6;
// bram[1943] = 10;
// bram[1944] = 16;
// bram[1945] = 23;
// bram[1946] = 32;
// bram[1947] = 41;
// bram[1948] = 51;
// bram[1949] = 62;
// bram[1950] = 73;
// bram[1951] = 85;
// bram[1952] = 98;
// bram[1953] = 111;
// bram[1954] = 124;
// bram[1955] = 137;
// bram[1956] = 150;
// bram[1957] = 163;
// bram[1958] = 175;
// bram[1959] = 187;
// bram[1960] = 198;
// bram[1961] = 208;
// bram[1962] = 218;
// bram[1963] = 226;
// bram[1964] = 234;
// bram[1965] = 240;
// bram[1966] = 246;
// bram[1967] = 249;
// bram[1968] = 252;
// bram[1969] = 253;
// bram[1970] = 253;
// bram[1971] = 252;
// bram[1972] = 249;
// bram[1973] = 245;
// bram[1974] = 240;
// bram[1975] = 233;
// bram[1976] = 226;
// bram[1977] = 217;
// bram[1978] = 208;
// bram[1979] = 197;
// bram[1980] = 186;
// bram[1981] = 174;
// bram[1982] = 162;
// bram[1983] = 149;
// bram[1984] = 136;
// bram[1985] = 123;
// bram[1986] = 110;
// bram[1987] = 97;
// bram[1988] = 85;
// bram[1989] = 73;
// bram[1990] = 61;
// bram[1991] = 50;
// bram[1992] = 40;
// bram[1993] = 31;
// bram[1994] = 23;
// bram[1995] = 16;
// bram[1996] = 10;
// bram[1997] = 6;
// bram[1998] = 2;
// bram[1999] = 0;
// bram[2000] = 0;
// bram[2001] = 0;
// bram[2002] = 2;
// bram[2003] = 6;
// bram[2004] = 10;
// bram[2005] = 16;
// bram[2006] = 23;
// bram[2007] = 31;
// bram[2008] = 40;
// bram[2009] = 50;
// bram[2010] = 61;
// bram[2011] = 73;
// bram[2012] = 85;
// bram[2013] = 97;
// bram[2014] = 110;
// bram[2015] = 123;
// bram[2016] = 136;
// bram[2017] = 149;
// bram[2018] = 162;
// bram[2019] = 174;
// bram[2020] = 186;
// bram[2021] = 197;
// bram[2022] = 208;
// bram[2023] = 217;
// bram[2024] = 226;
// bram[2025] = 233;
// bram[2026] = 240;
// bram[2027] = 245;
// bram[2028] = 249;
// bram[2029] = 252;
// bram[2030] = 253;
// bram[2031] = 253;
// bram[2032] = 252;
// bram[2033] = 249;
// bram[2034] = 246;
// bram[2035] = 240;
// bram[2036] = 234;
// bram[2037] = 226;
// bram[2038] = 218;
// bram[2039] = 208;
// bram[2040] = 198;
// bram[2041] = 187;
// bram[2042] = 175;
// bram[2043] = 163;
// bram[2044] = 150;
// bram[2045] = 137;
// bram[2046] = 124;
// bram[2047] = 111;
// bram[2048] = 98;
// bram[2049] = 85;
// bram[2050] = 73;
// bram[2051] = 62;
// bram[2052] = 51;
// bram[2053] = 41;
// bram[2054] = 32;
// bram[2055] = 23;
// bram[2056] = 16;
// bram[2057] = 10;
// bram[2058] = 6;
// bram[2059] = 2;
// bram[2060] = 0;
// bram[2061] = 0;
// bram[2062] = 0;
// bram[2063] = 2;
// bram[2064] = 5;
// bram[2065] = 10;
// bram[2066] = 15;
// bram[2067] = 22;
// bram[2068] = 30;
// bram[2069] = 39;
// bram[2070] = 49;
// bram[2071] = 60;
// bram[2072] = 72;
// bram[2073] = 84;
// bram[2074] = 96;
// bram[2075] = 109;
// bram[2076] = 122;
// bram[2077] = 135;
// bram[2078] = 148;
// bram[2079] = 161;
// bram[2080] = 173;
// bram[2081] = 185;
// bram[2082] = 196;
// bram[2083] = 207;
// bram[2084] = 217;
// bram[2085] = 225;
// bram[2086] = 233;
// bram[2087] = 240;
// bram[2088] = 245;
// bram[2089] = 249;
// bram[2090] = 252;
// bram[2091] = 253;
// bram[2092] = 253;
// bram[2093] = 252;
// bram[2094] = 250;
// bram[2095] = 246;
// bram[2096] = 241;
// bram[2097] = 234;
// bram[2098] = 227;
// bram[2099] = 218;
// bram[2100] = 209;
// bram[2101] = 199;
// bram[2102] = 188;
// bram[2103] = 176;
// bram[2104] = 163;
// bram[2105] = 151;
// bram[2106] = 138;
// bram[2107] = 125;
// bram[2108] = 112;
// bram[2109] = 99;
// bram[2110] = 86;
// bram[2111] = 74;
// bram[2112] = 63;
// bram[2113] = 52;
// bram[2114] = 41;
// bram[2115] = 32;
// bram[2116] = 24;
// bram[2117] = 17;
// bram[2118] = 11;
// bram[2119] = 6;
// bram[2120] = 3;
// bram[2121] = 0;
// bram[2122] = 0;
// bram[2123] = 0;
// bram[2124] = 2;
// bram[2125] = 5;
// bram[2126] = 9;
// bram[2127] = 15;
// bram[2128] = 22;
// bram[2129] = 30;
// bram[2130] = 39;
// bram[2131] = 49;
// bram[2132] = 59;
// bram[2133] = 71;
// bram[2134] = 83;
// bram[2135] = 95;
// bram[2136] = 108;
// bram[2137] = 121;
// bram[2138] = 134;
// bram[2139] = 147;
// bram[2140] = 160;
// bram[2141] = 172;
// bram[2142] = 184;
// bram[2143] = 196;
// bram[2144] = 206;
// bram[2145] = 216;
// bram[2146] = 225;
// bram[2147] = 232;
// bram[2148] = 239;
// bram[2149] = 245;
// bram[2150] = 249;
// bram[2151] = 252;
// bram[2152] = 253;
// bram[2153] = 253;
// bram[2154] = 252;
// bram[2155] = 250;
// bram[2156] = 246;
// bram[2157] = 241;
// bram[2158] = 235;
// bram[2159] = 228;
// bram[2160] = 219;
// bram[2161] = 210;
// bram[2162] = 199;
// bram[2163] = 188;
// bram[2164] = 177;
// bram[2165] = 164;
// bram[2166] = 152;
// bram[2167] = 139;
// bram[2168] = 126;
// bram[2169] = 113;
// bram[2170] = 100;
// bram[2171] = 87;
// bram[2172] = 75;
// bram[2173] = 63;
// bram[2174] = 52;
// bram[2175] = 42;
// bram[2176] = 33;
// bram[2177] = 25;
// bram[2178] = 17;
// bram[2179] = 11;
// bram[2180] = 6;
// bram[2181] = 3;
// bram[2182] = 0;
// bram[2183] = 0;
// bram[2184] = 0;
// bram[2185] = 2;
// bram[2186] = 5;
// bram[2187] = 9;
// bram[2188] = 15;
// bram[2189] = 21;
// bram[2190] = 29;
// bram[2191] = 38;
// bram[2192] = 48;
// bram[2193] = 59;
// bram[2194] = 70;
// bram[2195] = 82;
// bram[2196] = 95;
// bram[2197] = 107;
// bram[2198] = 120;
// bram[2199] = 133;
// bram[2200] = 146;
// bram[2201] = 159;
// bram[2202] = 172;
// bram[2203] = 184;
// bram[2204] = 195;
// bram[2205] = 206;
// bram[2206] = 215;
// bram[2207] = 224;
// bram[2208] = 232;
// bram[2209] = 239;
// bram[2210] = 244;
// bram[2211] = 248;
// bram[2212] = 251;
// bram[2213] = 253;
// bram[2214] = 253;
// bram[2215] = 252;
// bram[2216] = 250;
// bram[2217] = 246;
// bram[2218] = 241;
// bram[2219] = 235;
// bram[2220] = 228;
// bram[2221] = 220;
// bram[2222] = 210;
// bram[2223] = 200;
// bram[2224] = 189;
// bram[2225] = 177;
// bram[2226] = 165;
// bram[2227] = 153;
// bram[2228] = 140;
// bram[2229] = 127;
// bram[2230] = 114;
// bram[2231] = 101;
// bram[2232] = 88;
// bram[2233] = 76;
// bram[2234] = 64;
// bram[2235] = 53;
// bram[2236] = 43;
// bram[2237] = 33;
// bram[2238] = 25;
// bram[2239] = 18;
// bram[2240] = 12;
// bram[2241] = 7;
// bram[2242] = 3;
// bram[2243] = 1;
// bram[2244] = 0;
// bram[2245] = 0;
// bram[2246] = 1;
// bram[2247] = 4;
// bram[2248] = 9;
// bram[2249] = 14;
// bram[2250] = 21;
// bram[2251] = 29;
// bram[2252] = 38;
// bram[2253] = 47;
// bram[2254] = 58;
// bram[2255] = 69;
// bram[2256] = 81;
// bram[2257] = 94;
// bram[2258] = 106;
// bram[2259] = 119;
// bram[2260] = 132;
// bram[2261] = 145;
// bram[2262] = 158;
// bram[2263] = 171;
// bram[2264] = 183;
// bram[2265] = 194;
// bram[2266] = 205;
// bram[2267] = 215;
// bram[2268] = 224;
// bram[2269] = 231;
// bram[2270] = 238;
// bram[2271] = 244;
// bram[2272] = 248;
// bram[2273] = 251;
// bram[2274] = 253;
// bram[2275] = 253;
// bram[2276] = 253;
// bram[2277] = 250;
// bram[2278] = 247;
// bram[2279] = 242;
// bram[2280] = 236;
// bram[2281] = 229;
// bram[2282] = 220;
// bram[2283] = 211;
// bram[2284] = 201;
// bram[2285] = 190;
// bram[2286] = 178;
// bram[2287] = 166;
// bram[2288] = 153;
// bram[2289] = 141;
// bram[2290] = 127;
// bram[2291] = 114;
// bram[2292] = 102;
// bram[2293] = 89;
// bram[2294] = 77;
// bram[2295] = 65;
// bram[2296] = 54;
// bram[2297] = 43;
// bram[2298] = 34;
// bram[2299] = 26;
// bram[2300] = 18;
// bram[2301] = 12;
// bram[2302] = 7;
// bram[2303] = 3;
// bram[2304] = 1;
// bram[2305] = 0;
// bram[2306] = 0;
// bram[2307] = 1;
// bram[2308] = 4;
// bram[2309] = 8;
// bram[2310] = 14;
// bram[2311] = 20;
// bram[2312] = 28;
// bram[2313] = 37;
// bram[2314] = 47;
// bram[2315] = 57;
// bram[2316] = 68;
// bram[2317] = 80;
// bram[2318] = 93;
// bram[2319] = 106;
// bram[2320] = 119;
// bram[2321] = 132;
// bram[2322] = 145;
// bram[2323] = 157;
// bram[2324] = 170;
// bram[2325] = 182;
// bram[2326] = 193;
// bram[2327] = 204;
// bram[2328] = 214;
// bram[2329] = 223;
// bram[2330] = 231;
// bram[2331] = 238;
// bram[2332] = 244;
// bram[2333] = 248;
// bram[2334] = 251;
// bram[2335] = 253;
// bram[2336] = 253;
// bram[2337] = 253;
// bram[2338] = 250;
// bram[2339] = 247;
// bram[2340] = 242;
// bram[2341] = 236;
// bram[2342] = 229;
// bram[2343] = 221;
// bram[2344] = 212;
// bram[2345] = 202;
// bram[2346] = 191;
// bram[2347] = 179;
// bram[2348] = 167;
// bram[2349] = 154;
// bram[2350] = 141;
// bram[2351] = 128;
// bram[2352] = 115;
// bram[2353] = 102;
// bram[2354] = 90;
// bram[2355] = 77;
// bram[2356] = 66;
// bram[2357] = 55;
// bram[2358] = 44;
// bram[2359] = 35;
// bram[2360] = 26;
// bram[2361] = 19;
// bram[2362] = 12;
// bram[2363] = 7;
// bram[2364] = 3;
// bram[2365] = 1;
// bram[2366] = 0;
// bram[2367] = 0;
// bram[2368] = 1;
// bram[2369] = 4;
// bram[2370] = 8;
// bram[2371] = 13;
// bram[2372] = 20;
// bram[2373] = 28;
// bram[2374] = 36;
// bram[2375] = 46;
// bram[2376] = 56;
// bram[2377] = 68;
// bram[2378] = 80;
// bram[2379] = 92;
// bram[2380] = 105;
// bram[2381] = 118;
// bram[2382] = 131;
// bram[2383] = 144;
// bram[2384] = 157;
// bram[2385] = 169;
// bram[2386] = 181;
// bram[2387] = 193;
// bram[2388] = 203;
// bram[2389] = 213;
// bram[2390] = 222;
// bram[2391] = 230;
// bram[2392] = 237;
// bram[2393] = 243;
// bram[2394] = 248;
// bram[2395] = 251;
// bram[2396] = 253;
// bram[2397] = 253;
// bram[2398] = 253;
// bram[2399] = 251;
// bram[2400] = 247;
// bram[2401] = 243;
// bram[2402] = 237;
// bram[2403] = 230;
// bram[2404] = 221;
// bram[2405] = 212;
// bram[2406] = 202;
// bram[2407] = 191;
// bram[2408] = 180;
// bram[2409] = 168;
// bram[2410] = 155;
// bram[2411] = 142;
// bram[2412] = 129;
// bram[2413] = 116;
// bram[2414] = 103;
// bram[2415] = 91;
// bram[2416] = 78;
// bram[2417] = 66;
// bram[2418] = 55;
// bram[2419] = 45;
// bram[2420] = 35;
// bram[2421] = 27;
// bram[2422] = 19;
// bram[2423] = 13;
// bram[2424] = 8;
// bram[2425] = 4;
// bram[2426] = 1;
// bram[2427] = 0;
// bram[2428] = 0;
// bram[2429] = 1;
// bram[2430] = 4;
// bram[2431] = 8;
// bram[2432] = 13;
// bram[2433] = 19;
// bram[2434] = 27;
// bram[2435] = 36;
// bram[2436] = 45;
// bram[2437] = 56;
// bram[2438] = 67;
// bram[2439] = 79;
// bram[2440] = 91;
// bram[2441] = 104;
// bram[2442] = 117;
// bram[2443] = 130;
// bram[2444] = 143;
// bram[2445] = 156;
// bram[2446] = 168;
// bram[2447] = 180;
// bram[2448] = 192;
// bram[2449] = 203;
// bram[2450] = 213;
// bram[2451] = 222;
// bram[2452] = 230;
// bram[2453] = 237;
// bram[2454] = 243;
// bram[2455] = 247;
// bram[2456] = 251;
// bram[2457] = 253;
// bram[2458] = 253;
// bram[2459] = 253;
// bram[2460] = 251;
// bram[2461] = 248;
// bram[2462] = 243;
// bram[2463] = 237;
// bram[2464] = 230;
// bram[2465] = 222;
// bram[2466] = 213;
// bram[2467] = 203;
// bram[2468] = 192;
// bram[2469] = 181;
// bram[2470] = 169;
// bram[2471] = 156;
// bram[2472] = 143;
// bram[2473] = 130;
// bram[2474] = 117;
// bram[2475] = 104;
// bram[2476] = 91;
// bram[2477] = 79;
// bram[2478] = 67;
// bram[2479] = 56;
// bram[2480] = 46;
// bram[2481] = 36;
// bram[2482] = 27;
// bram[2483] = 20;
// bram[2484] = 13;
// bram[2485] = 8;
// bram[2486] = 4;
// bram[2487] = 1;
// bram[2488] = 0;
// bram[2489] = 0;
// bram[2490] = 1;
// bram[2491] = 4;
// bram[2492] = 7;
// bram[2493] = 13;
// bram[2494] = 19;
// bram[2495] = 26;
// bram[2496] = 35;
// bram[2497] = 45;
// bram[2498] = 55;
// bram[2499] = 66;
// bram[2500] = 78;
// bram[2501] = 90;
// bram[2502] = 103;
// bram[2503] = 116;
// bram[2504] = 129;
// bram[2505] = 142;
// bram[2506] = 155;
// bram[2507] = 167;
// bram[2508] = 179;
// bram[2509] = 191;
// bram[2510] = 202;
// bram[2511] = 212;
// bram[2512] = 221;
// bram[2513] = 229;
// bram[2514] = 237;
// bram[2515] = 242;
// bram[2516] = 247;
// bram[2517] = 251;
// bram[2518] = 253;
// bram[2519] = 253;
// bram[2520] = 253;
// bram[2521] = 251;
// bram[2522] = 248;
// bram[2523] = 243;
// bram[2524] = 238;
// bram[2525] = 231;
// bram[2526] = 223;
// bram[2527] = 214;
// bram[2528] = 204;
// bram[2529] = 193;
// bram[2530] = 181;
// bram[2531] = 169;
// bram[2532] = 157;
// bram[2533] = 144;
// bram[2534] = 131;
// bram[2535] = 118;
// bram[2536] = 105;
// bram[2537] = 92;
// bram[2538] = 80;
// bram[2539] = 68;
// bram[2540] = 57;
// bram[2541] = 46;
// bram[2542] = 37;
// bram[2543] = 28;
// bram[2544] = 20;
// bram[2545] = 14;
// bram[2546] = 8;
// bram[2547] = 4;
// bram[2548] = 1;
// bram[2549] = 0;
// bram[2550] = 0;
// bram[2551] = 1;
// bram[2552] = 3;
// bram[2553] = 7;
// bram[2554] = 12;
// bram[2555] = 18;
// bram[2556] = 26;
// bram[2557] = 34;
// bram[2558] = 44;
// bram[2559] = 54;
// bram[2560] = 65;
// bram[2561] = 77;
// bram[2562] = 89;
// bram[2563] = 102;
// bram[2564] = 115;
// bram[2565] = 128;
// bram[2566] = 141;
// bram[2567] = 154;
// bram[2568] = 167;
// bram[2569] = 179;
// bram[2570] = 190;
// bram[2571] = 201;
// bram[2572] = 211;
// bram[2573] = 221;
// bram[2574] = 229;
// bram[2575] = 236;
// bram[2576] = 242;
// bram[2577] = 247;
// bram[2578] = 250;
// bram[2579] = 253;
// bram[2580] = 253;
// bram[2581] = 253;
// bram[2582] = 251;
// bram[2583] = 248;
// bram[2584] = 244;
// bram[2585] = 238;
// bram[2586] = 231;
// bram[2587] = 223;
// bram[2588] = 214;
// bram[2589] = 204;
// bram[2590] = 194;
// bram[2591] = 182;
// bram[2592] = 170;
// bram[2593] = 158;
// bram[2594] = 145;
// bram[2595] = 132;
// bram[2596] = 119;
// bram[2597] = 106;
// bram[2598] = 93;
// bram[2599] = 81;
// bram[2600] = 69;
// bram[2601] = 58;
// bram[2602] = 47;
// bram[2603] = 37;
// bram[2604] = 28;
// bram[2605] = 21;
// bram[2606] = 14;
// bram[2607] = 9;
// bram[2608] = 4;
// bram[2609] = 1;
// bram[2610] = 0;
// bram[2611] = 0;
// bram[2612] = 1;
// bram[2613] = 3;
// bram[2614] = 7;
// bram[2615] = 12;
// bram[2616] = 18;
// bram[2617] = 25;
// bram[2618] = 34;
// bram[2619] = 43;
// bram[2620] = 53;
// bram[2621] = 65;
// bram[2622] = 76;
// bram[2623] = 88;
// bram[2624] = 101;
// bram[2625] = 114;
// bram[2626] = 127;
// bram[2627] = 140;
// bram[2628] = 153;
// bram[2629] = 166;
// bram[2630] = 178;
// bram[2631] = 190;
// bram[2632] = 201;
// bram[2633] = 211;
// bram[2634] = 220;
// bram[2635] = 228;
// bram[2636] = 236;
// bram[2637] = 242;
// bram[2638] = 247;
// bram[2639] = 250;
// bram[2640] = 252;
// bram[2641] = 253;
// bram[2642] = 253;
// bram[2643] = 251;
// bram[2644] = 248;
// bram[2645] = 244;
// bram[2646] = 238;
// bram[2647] = 232;
// bram[2648] = 224;
// bram[2649] = 215;
// bram[2650] = 205;
// bram[2651] = 194;
// bram[2652] = 183;
// bram[2653] = 171;
// bram[2654] = 159;
// bram[2655] = 146;
// bram[2656] = 133;
// bram[2657] = 120;
// bram[2658] = 107;
// bram[2659] = 94;
// bram[2660] = 82;
// bram[2661] = 70;
// bram[2662] = 58;
// bram[2663] = 48;
// bram[2664] = 38;
// bram[2665] = 29;
// bram[2666] = 21;
// bram[2667] = 14;
// bram[2668] = 9;
// bram[2669] = 5;
// bram[2670] = 2;
// bram[2671] = 0;
// bram[2672] = 0;
// bram[2673] = 1;
// bram[2674] = 3;
// bram[2675] = 7;
// bram[2676] = 11;
// bram[2677] = 18;
// bram[2678] = 25;
// bram[2679] = 33;
// bram[2680] = 43;
// bram[2681] = 53;
// bram[2682] = 64;
// bram[2683] = 75;
// bram[2684] = 88;
// bram[2685] = 100;
// bram[2686] = 113;
// bram[2687] = 126;
// bram[2688] = 139;
// bram[2689] = 152;
// bram[2690] = 165;
// bram[2691] = 177;
// bram[2692] = 189;
// bram[2693] = 200;
// bram[2694] = 210;
// bram[2695] = 219;
// bram[2696] = 228;
// bram[2697] = 235;
// bram[2698] = 241;
// bram[2699] = 246;
// bram[2700] = 250;
// bram[2701] = 252;
// bram[2702] = 253;
// bram[2703] = 253;
// bram[2704] = 252;
// bram[2705] = 249;
// bram[2706] = 244;
// bram[2707] = 239;
// bram[2708] = 232;
// bram[2709] = 224;
// bram[2710] = 216;
// bram[2711] = 206;
// bram[2712] = 195;
// bram[2713] = 184;
// bram[2714] = 172;
// bram[2715] = 160;
// bram[2716] = 147;
// bram[2717] = 134;
// bram[2718] = 121;
// bram[2719] = 108;
// bram[2720] = 95;
// bram[2721] = 82;
// bram[2722] = 70;
// bram[2723] = 59;
// bram[2724] = 48;
// bram[2725] = 38;
// bram[2726] = 30;
// bram[2727] = 22;
// bram[2728] = 15;
// bram[2729] = 9;
// bram[2730] = 5;
// bram[2731] = 2;
// bram[2732] = 0;
// bram[2733] = 0;
// bram[2734] = 0;
// bram[2735] = 3;
// bram[2736] = 6;
// bram[2737] = 11;
// bram[2738] = 17;
// bram[2739] = 24;
// bram[2740] = 33;
// bram[2741] = 42;
// bram[2742] = 52;
// bram[2743] = 63;
// bram[2744] = 75;
// bram[2745] = 87;
// bram[2746] = 99;
// bram[2747] = 112;
// bram[2748] = 125;
// bram[2749] = 138;
// bram[2750] = 151;
// bram[2751] = 164;
// bram[2752] = 176;
// bram[2753] = 188;
// bram[2754] = 199;
// bram[2755] = 209;
// bram[2756] = 219;
// bram[2757] = 227;
// bram[2758] = 235;
// bram[2759] = 241;
// bram[2760] = 246;
// bram[2761] = 250;
// bram[2762] = 252;
// bram[2763] = 253;
// bram[2764] = 253;
// bram[2765] = 252;
// bram[2766] = 249;
// bram[2767] = 245;
// bram[2768] = 239;
// bram[2769] = 233;
// bram[2770] = 225;
// bram[2771] = 216;
// bram[2772] = 207;
// bram[2773] = 196;
// bram[2774] = 185;
// bram[2775] = 173;
// bram[2776] = 160;
// bram[2777] = 148;
// bram[2778] = 135;
// bram[2779] = 122;
// bram[2780] = 109;
// bram[2781] = 96;
// bram[2782] = 83;
// bram[2783] = 71;
// bram[2784] = 60;
// bram[2785] = 49;
// bram[2786] = 39;
// bram[2787] = 30;
// bram[2788] = 22;
// bram[2789] = 15;
// bram[2790] = 10;
// bram[2791] = 5;
// bram[2792] = 2;
// bram[2793] = 0;
// bram[2794] = 0;
// bram[2795] = 0;
// bram[2796] = 2;
// bram[2797] = 6;
// bram[2798] = 11;
// bram[2799] = 17;
// bram[2800] = 24;
// bram[2801] = 32;
// bram[2802] = 41;
// bram[2803] = 51;
// bram[2804] = 62;
// bram[2805] = 74;
// bram[2806] = 86;
// bram[2807] = 99;
// bram[2808] = 111;
// bram[2809] = 124;
// bram[2810] = 137;
// bram[2811] = 150;
// bram[2812] = 163;
// bram[2813] = 175;
// bram[2814] = 187;
// bram[2815] = 198;
// bram[2816] = 209;
// bram[2817] = 218;
// bram[2818] = 227;
// bram[2819] = 234;
// bram[2820] = 241;
// bram[2821] = 246;
// bram[2822] = 250;
// bram[2823] = 252;
// bram[2824] = 253;
// bram[2825] = 253;
// bram[2826] = 252;
// bram[2827] = 249;
// bram[2828] = 245;
// bram[2829] = 240;
// bram[2830] = 233;
// bram[2831] = 226;
// bram[2832] = 217;
// bram[2833] = 207;
// bram[2834] = 197;
// bram[2835] = 185;
// bram[2836] = 174;
// bram[2837] = 161;
// bram[2838] = 149;
// bram[2839] = 136;
// bram[2840] = 123;
// bram[2841] = 109;
// bram[2842] = 97;
// bram[2843] = 84;
// bram[2844] = 72;
// bram[2845] = 61;
// bram[2846] = 50;
// bram[2847] = 40;
// bram[2848] = 31;
// bram[2849] = 23;
// bram[2850] = 16;
// bram[2851] = 10;
// bram[2852] = 5;
// bram[2853] = 2;
// bram[2854] = 0;
// bram[2855] = 0;
// bram[2856] = 0;
// bram[2857] = 2;
// bram[2858] = 6;
// bram[2859] = 10;
// bram[2860] = 16;
// bram[2861] = 23;
// bram[2862] = 31;
// bram[2863] = 41;
// bram[2864] = 51;
// bram[2865] = 61;
// bram[2866] = 73;
// bram[2867] = 85;
// bram[2868] = 98;
// bram[2869] = 110;
// bram[2870] = 124;
// bram[2871] = 137;
// bram[2872] = 150;
// bram[2873] = 162;
// bram[2874] = 175;
// bram[2875] = 186;
// bram[2876] = 198;
// bram[2877] = 208;
// bram[2878] = 218;
// bram[2879] = 226;
// bram[2880] = 234;
// bram[2881] = 240;
// bram[2882] = 245;
// bram[2883] = 249;
// bram[2884] = 252;
// bram[2885] = 253;
// bram[2886] = 253;
// bram[2887] = 252;
// bram[2888] = 249;
// bram[2889] = 245;
// bram[2890] = 240;
// bram[2891] = 234;
// bram[2892] = 226;
// bram[2893] = 217;
// bram[2894] = 208;
// bram[2895] = 197;
// bram[2896] = 186;
// bram[2897] = 174;
// bram[2898] = 162;
// bram[2899] = 149;
// bram[2900] = 136;
// bram[2901] = 123;
// bram[2902] = 110;
// bram[2903] = 98;
// bram[2904] = 85;
// bram[2905] = 73;
// bram[2906] = 61;
// bram[2907] = 50;
// bram[2908] = 40;
// bram[2909] = 31;
// bram[2910] = 23;
// bram[2911] = 16;
// bram[2912] = 10;
// bram[2913] = 6;
// bram[2914] = 2;
// bram[2915] = 0;
// bram[2916] = 0;
// bram[2917] = 0;
// bram[2918] = 2;
// bram[2919] = 5;
// bram[2920] = 10;
// bram[2921] = 16;
// bram[2922] = 23;
// bram[2923] = 31;
// bram[2924] = 40;
// bram[2925] = 50;
// bram[2926] = 61;
// bram[2927] = 72;
// bram[2928] = 84;
// bram[2929] = 97;
// bram[2930] = 110;
// bram[2931] = 123;
// bram[2932] = 136;
// bram[2933] = 149;
// bram[2934] = 161;
// bram[2935] = 174;
// bram[2936] = 186;
// bram[2937] = 197;
// bram[2938] = 207;
// bram[2939] = 217;
// bram[2940] = 226;
// bram[2941] = 233;
// bram[2942] = 240;
// bram[2943] = 245;
// bram[2944] = 249;
// bram[2945] = 252;
// bram[2946] = 253;
// bram[2947] = 253;
// bram[2948] = 252;
// bram[2949] = 250;
// bram[2950] = 246;
// bram[2951] = 241;
// bram[2952] = 234;
// bram[2953] = 227;
// bram[2954] = 218;
// bram[2955] = 209;
// bram[2956] = 198;
// bram[2957] = 187;
// bram[2958] = 175;
// bram[2959] = 163;
// bram[2960] = 150;
// bram[2961] = 137;
// bram[2962] = 124;
// bram[2963] = 111;
// bram[2964] = 98;
// bram[2965] = 86;
// bram[2966] = 74;
// bram[2967] = 62;
// bram[2968] = 51;
// bram[2969] = 41;
// bram[2970] = 32;
// bram[2971] = 24;
// bram[2972] = 17;
// bram[2973] = 11;
// bram[2974] = 6;
// bram[2975] = 2;
// bram[2976] = 0;
// bram[2977] = 0;
// bram[2978] = 0;
// bram[2979] = 2;
// bram[2980] = 5;
// bram[2981] = 10;
// bram[2982] = 15;
// bram[2983] = 22;
// bram[2984] = 30;
// bram[2985] = 39;
// bram[2986] = 49;
// bram[2987] = 60;
// bram[2988] = 71;
// bram[2989] = 83;
// bram[2990] = 96;
// bram[2991] = 109;
// bram[2992] = 122;
// bram[2993] = 135;
// bram[2994] = 148;
// bram[2995] = 160;
// bram[2996] = 173;
// bram[2997] = 185;
// bram[2998] = 196;
// bram[2999] = 207;
// bram[3000] = 216;
// bram[3001] = 225;
// bram[3002] = 233;
// bram[3003] = 239;
// bram[3004] = 245;
// bram[3005] = 249;
// bram[3006] = 252;
// bram[3007] = 253;
// bram[3008] = 253;
// bram[3009] = 252;
// bram[3010] = 250;
// bram[3011] = 246;
// bram[3012] = 241;
// bram[3013] = 235;
// bram[3014] = 227;
// bram[3015] = 219;
// bram[3016] = 209;
// bram[3017] = 199;
// bram[3018] = 188;
// bram[3019] = 176;
// bram[3020] = 164;
// bram[3021] = 151;
// bram[3022] = 138;
// bram[3023] = 125;
// bram[3024] = 112;
// bram[3025] = 99;
// bram[3026] = 87;
// bram[3027] = 75;
// bram[3028] = 63;
// bram[3029] = 52;
// bram[3030] = 42;
// bram[3031] = 32;
// bram[3032] = 24;
// bram[3033] = 17;
// bram[3034] = 11;
// bram[3035] = 6;
// bram[3036] = 3;
// bram[3037] = 0;
// bram[3038] = 0;
// bram[3039] = 0;
// bram[3040] = 2;
// bram[3041] = 5;
// bram[3042] = 9;
// bram[3043] = 15;
// bram[3044] = 22;
// bram[3045] = 30;
// bram[3046] = 39;
// bram[3047] = 48;
// bram[3048] = 59;
// bram[3049] = 71;
// bram[3050] = 83;
// bram[3051] = 95;
// bram[3052] = 108;
// bram[3053] = 121;
// bram[3054] = 134;
// bram[3055] = 147;
// bram[3056] = 160;
// bram[3057] = 172;
// bram[3058] = 184;
// bram[3059] = 195;
// bram[3060] = 206;
// bram[3061] = 216;
// bram[3062] = 224;
// bram[3063] = 232;
// bram[3064] = 239;
// bram[3065] = 244;
// bram[3066] = 249;
// bram[3067] = 252;
// bram[3068] = 253;
// bram[3069] = 253;
// bram[3070] = 252;
// bram[3071] = 250;
// bram[3072] = 246;
// bram[3073] = 241;
// bram[3074] = 235;
// bram[3075] = 228;
// bram[3076] = 219;
// bram[3077] = 210;
// bram[3078] = 200;
// bram[3079] = 189;
// bram[3080] = 177;
// bram[3081] = 165;
// bram[3082] = 152;
// bram[3083] = 139;
// bram[3084] = 126;
// bram[3085] = 113;
// bram[3086] = 100;
// bram[3087] = 88;
// bram[3088] = 75;
// bram[3089] = 64;
// bram[3090] = 53;
// bram[3091] = 42;
// bram[3092] = 33;
// bram[3093] = 25;
// bram[3094] = 17;
// bram[3095] = 11;
// bram[3096] = 6;
// bram[3097] = 3;
// bram[3098] = 1;
// bram[3099] = 0;
// bram[3100] = 0;
// bram[3101] = 2;
// bram[3102] = 5;
// bram[3103] = 9;
// bram[3104] = 14;
// bram[3105] = 21;
// bram[3106] = 29;
// bram[3107] = 38;
// bram[3108] = 48;
// bram[3109] = 58;
// bram[3110] = 70;
// bram[3111] = 82;
// bram[3112] = 94;
// bram[3113] = 107;
// bram[3114] = 120;
// bram[3115] = 133;
// bram[3116] = 146;
// bram[3117] = 159;
// bram[3118] = 171;
// bram[3119] = 183;
// bram[3120] = 195;
// bram[3121] = 205;
// bram[3122] = 215;
// bram[3123] = 224;
// bram[3124] = 232;
// bram[3125] = 239;
// bram[3126] = 244;
// bram[3127] = 248;
// bram[3128] = 251;
// bram[3129] = 253;
// bram[3130] = 253;
// bram[3131] = 252;
// bram[3132] = 250;
// bram[3133] = 247;
// bram[3134] = 242;
// bram[3135] = 236;
// bram[3136] = 228;
// bram[3137] = 220;
// bram[3138] = 211;
// bram[3139] = 200;
// bram[3140] = 189;
// bram[3141] = 178;
// bram[3142] = 166;
// bram[3143] = 153;
// bram[3144] = 140;
// bram[3145] = 127;
// bram[3146] = 114;
// bram[3147] = 101;
// bram[3148] = 88;
// bram[3149] = 76;
// bram[3150] = 64;
// bram[3151] = 53;
// bram[3152] = 43;
// bram[3153] = 34;
// bram[3154] = 25;
// bram[3155] = 18;
// bram[3156] = 12;
// bram[3157] = 7;
// bram[3158] = 3;
// bram[3159] = 1;
// bram[3160] = 0;
// bram[3161] = 0;
// bram[3162] = 1;
// bram[3163] = 4;
// bram[3164] = 9;
// bram[3165] = 14;
// bram[3166] = 21;
// bram[3167] = 28;
// bram[3168] = 37;
// bram[3169] = 47;
// bram[3170] = 58;
// bram[3171] = 69;
// bram[3172] = 81;
// bram[3173] = 93;
// bram[3174] = 106;
// bram[3175] = 119;
// bram[3176] = 132;
// bram[3177] = 145;
// bram[3178] = 158;
// bram[3179] = 170;
// bram[3180] = 182;
// bram[3181] = 194;
// bram[3182] = 204;
// bram[3183] = 214;
// bram[3184] = 223;
// bram[3185] = 231;
// bram[3186] = 238;
// bram[3187] = 244;
// bram[3188] = 248;
// bram[3189] = 251;
// bram[3190] = 253;
// bram[3191] = 253;
// bram[3192] = 253;
// bram[3193] = 250;
// bram[3194] = 247;
// bram[3195] = 242;
// bram[3196] = 236;
// bram[3197] = 229;
// bram[3198] = 221;
// bram[3199] = 211;
// bram[3200] = 201;
// bram[3201] = 190;
// bram[3202] = 179;
// bram[3203] = 166;
// bram[3204] = 154;
// bram[3205] = 141;
// bram[3206] = 128;
// bram[3207] = 115;
// bram[3208] = 102;
// bram[3209] = 89;
// bram[3210] = 77;
// bram[3211] = 65;
// bram[3212] = 54;
// bram[3213] = 44;
// bram[3214] = 34;
// bram[3215] = 26;
// bram[3216] = 18;
// bram[3217] = 12;
// bram[3218] = 7;
// bram[3219] = 3;
// bram[3220] = 1;
// bram[3221] = 0;
// bram[3222] = 0;
// bram[3223] = 1;
// bram[3224] = 4;
// bram[3225] = 8;
// bram[3226] = 14;
// bram[3227] = 20;
// bram[3228] = 28;
// bram[3229] = 37;
// bram[3230] = 46;
// bram[3231] = 57;
// bram[3232] = 68;
// bram[3233] = 80;
// bram[3234] = 92;
// bram[3235] = 105;
// bram[3236] = 118;
// bram[3237] = 131;
// bram[3238] = 144;
// bram[3239] = 157;
// bram[3240] = 170;
// bram[3241] = 182;
// bram[3242] = 193;
// bram[3243] = 204;
// bram[3244] = 214;
// bram[3245] = 223;
// bram[3246] = 231;
// bram[3247] = 238;
// bram[3248] = 243;
// bram[3249] = 248;
// bram[3250] = 251;
// bram[3251] = 253;
// bram[3252] = 253;
// bram[3253] = 253;
// bram[3254] = 251;
// bram[3255] = 247;
// bram[3256] = 242;
// bram[3257] = 236;
// bram[3258] = 229;
// bram[3259] = 221;
// bram[3260] = 212;
// bram[3261] = 202;
// bram[3262] = 191;
// bram[3263] = 179;
// bram[3264] = 167;
// bram[3265] = 155;
// bram[3266] = 142;
// bram[3267] = 129;
// bram[3268] = 116;
// bram[3269] = 103;
// bram[3270] = 90;
// bram[3271] = 78;
// bram[3272] = 66;
// bram[3273] = 55;
// bram[3274] = 44;
// bram[3275] = 35;
// bram[3276] = 26;
// bram[3277] = 19;
// bram[3278] = 13;
// bram[3279] = 7;
// bram[3280] = 3;
// bram[3281] = 1;
// bram[3282] = 0;
// bram[3283] = 0;
// bram[3284] = 1;
// bram[3285] = 4;
// bram[3286] = 8;
// bram[3287] = 13;
// bram[3288] = 20;
// bram[3289] = 27;
// bram[3290] = 36;
// bram[3291] = 46;
// bram[3292] = 56;
// bram[3293] = 67;
// bram[3294] = 79;
// bram[3295] = 92;
// bram[3296] = 104;
// bram[3297] = 117;
// bram[3298] = 130;
// bram[3299] = 143;
// bram[3300] = 156;
// bram[3301] = 169;
// bram[3302] = 181;
// bram[3303] = 192;
// bram[3304] = 203;
// bram[3305] = 213;
// bram[3306] = 222;
// bram[3307] = 230;
// bram[3308] = 237;
// bram[3309] = 243;
// bram[3310] = 248;
// bram[3311] = 251;
// bram[3312] = 253;
// bram[3313] = 253;
// bram[3314] = 253;
// bram[3315] = 251;
// bram[3316] = 247;
// bram[3317] = 243;
// bram[3318] = 237;
// bram[3319] = 230;
// bram[3320] = 222;
// bram[3321] = 213;
// bram[3322] = 203;
// bram[3323] = 192;
// bram[3324] = 180;
// bram[3325] = 168;
// bram[3326] = 156;
// bram[3327] = 143;
// bram[3328] = 130;
// bram[3329] = 117;
// bram[3330] = 104;
// bram[3331] = 91;
// bram[3332] = 79;
// bram[3333] = 67;
// bram[3334] = 56;
// bram[3335] = 45;
// bram[3336] = 36;
// bram[3337] = 27;
// bram[3338] = 19;
// bram[3339] = 13;
// bram[3340] = 8;
// bram[3341] = 4;
// bram[3342] = 1;
// bram[3343] = 0;
// bram[3344] = 0;
// bram[3345] = 1;
// bram[3346] = 4;
// bram[3347] = 8;
// bram[3348] = 13;
// bram[3349] = 19;
// bram[3350] = 27;
// bram[3351] = 35;
// bram[3352] = 45;
// bram[3353] = 55;
// bram[3354] = 67;
// bram[3355] = 78;
// bram[3356] = 91;
// bram[3357] = 103;
// bram[3358] = 116;
// bram[3359] = 129;
// bram[3360] = 142;
// bram[3361] = 155;
// bram[3362] = 168;
// bram[3363] = 180;
// bram[3364] = 191;
// bram[3365] = 202;
// bram[3366] = 212;
// bram[3367] = 222;
// bram[3368] = 230;
// bram[3369] = 237;
// bram[3370] = 243;
// bram[3371] = 247;
// bram[3372] = 251;
// bram[3373] = 253;
// bram[3374] = 253;
// bram[3375] = 253;
// bram[3376] = 251;
// bram[3377] = 248;
// bram[3378] = 243;
// bram[3379] = 237;
// bram[3380] = 230;
// bram[3381] = 222;
// bram[3382] = 213;
// bram[3383] = 203;
// bram[3384] = 193;
// bram[3385] = 181;
// bram[3386] = 169;
// bram[3387] = 156;
// bram[3388] = 144;
// bram[3389] = 131;
// bram[3390] = 118;
// bram[3391] = 105;
// bram[3392] = 92;
// bram[3393] = 79;
// bram[3394] = 68;
// bram[3395] = 56;
// bram[3396] = 46;
// bram[3397] = 36;
// bram[3398] = 28;
// bram[3399] = 20;
// bram[3400] = 13;
// bram[3401] = 8;
// bram[3402] = 4;
// bram[3403] = 1;
// bram[3404] = 0;
// bram[3405] = 0;
// bram[3406] = 1;
// bram[3407] = 3;
// bram[3408] = 7;
// bram[3409] = 12;
// bram[3410] = 19;
// bram[3411] = 26;
// bram[3412] = 35;
// bram[3413] = 44;
// bram[3414] = 55;
// bram[3415] = 66;
// bram[3416] = 78;
// bram[3417] = 90;
// bram[3418] = 103;
// bram[3419] = 115;
// bram[3420] = 128;
// bram[3421] = 142;
// bram[3422] = 154;
// bram[3423] = 167;
// bram[3424] = 179;
// bram[3425] = 191;
// bram[3426] = 202;
// bram[3427] = 212;
// bram[3428] = 221;
// bram[3429] = 229;
// bram[3430] = 236;
// bram[3431] = 242;
// bram[3432] = 247;
// bram[3433] = 251;
// bram[3434] = 253;
// bram[3435] = 253;
// bram[3436] = 253;
// bram[3437] = 251;
// bram[3438] = 248;
// bram[3439] = 243;
// bram[3440] = 238;
// bram[3441] = 231;
// bram[3442] = 223;
// bram[3443] = 214;
// bram[3444] = 204;
// bram[3445] = 193;
// bram[3446] = 182;
// bram[3447] = 170;
// bram[3448] = 157;
// bram[3449] = 144;
// bram[3450] = 131;
// bram[3451] = 118;
// bram[3452] = 105;
// bram[3453] = 93;
// bram[3454] = 80;
// bram[3455] = 68;
// bram[3456] = 57;
// bram[3457] = 47;
// bram[3458] = 37;
// bram[3459] = 28;
// bram[3460] = 20;
// bram[3461] = 14;
// bram[3462] = 8;
// bram[3463] = 4;
// bram[3464] = 1;
// bram[3465] = 0;
// bram[3466] = 0;
// bram[3467] = 1;
// bram[3468] = 3;
// bram[3469] = 7;
// bram[3470] = 12;
// bram[3471] = 18;
// bram[3472] = 26;
// bram[3473] = 34;
// bram[3474] = 44;
// bram[3475] = 54;
// bram[3476] = 65;
// bram[3477] = 77;
// bram[3478] = 89;
// bram[3479] = 102;
// bram[3480] = 115;
// bram[3481] = 128;
// bram[3482] = 141;
// bram[3483] = 154;
// bram[3484] = 166;
// bram[3485] = 178;
// bram[3486] = 190;
// bram[3487] = 201;
// bram[3488] = 211;
// bram[3489] = 220;
// bram[3490] = 229;
// bram[3491] = 236;
// bram[3492] = 242;
// bram[3493] = 247;
// bram[3494] = 250;
// bram[3495] = 253;
// bram[3496] = 253;
// bram[3497] = 253;
// bram[3498] = 251;
// bram[3499] = 248;
// bram[3500] = 244;
// bram[3501] = 238;
// bram[3502] = 231;
// bram[3503] = 224;
// bram[3504] = 215;
// bram[3505] = 205;
// bram[3506] = 194;
// bram[3507] = 183;
// bram[3508] = 171;
// bram[3509] = 158;
// bram[3510] = 145;
// bram[3511] = 132;
// bram[3512] = 119;
// bram[3513] = 106;
// bram[3514] = 94;
// bram[3515] = 81;
// bram[3516] = 69;
// bram[3517] = 58;
// bram[3518] = 47;
// bram[3519] = 37;
// bram[3520] = 29;
// bram[3521] = 21;
// bram[3522] = 14;
// bram[3523] = 9;
// bram[3524] = 4;
// bram[3525] = 1;
// bram[3526] = 0;
// bram[3527] = 0;
// bram[3528] = 1;
// bram[3529] = 3;
// bram[3530] = 7;
// bram[3531] = 12;
// bram[3532] = 18;
// bram[3533] = 25;
// bram[3534] = 34;
// bram[3535] = 43;
// bram[3536] = 53;
// bram[3537] = 64;
// bram[3538] = 76;
// bram[3539] = 88;
// bram[3540] = 101;
// bram[3541] = 114;
// bram[3542] = 127;
// bram[3543] = 140;
// bram[3544] = 153;
// bram[3545] = 165;
// bram[3546] = 177;
// bram[3547] = 189;
// bram[3548] = 200;
// bram[3549] = 210;
// bram[3550] = 220;
// bram[3551] = 228;
// bram[3552] = 235;
// bram[3553] = 242;
// bram[3554] = 246;
// bram[3555] = 250;
// bram[3556] = 252;
// bram[3557] = 253;
// bram[3558] = 253;
// bram[3559] = 251;
// bram[3560] = 248;
// bram[3561] = 244;
// bram[3562] = 239;
// bram[3563] = 232;
// bram[3564] = 224;
// bram[3565] = 215;
// bram[3566] = 205;
// bram[3567] = 195;
// bram[3568] = 183;
// bram[3569] = 171;
// bram[3570] = 159;
// bram[3571] = 146;
// bram[3572] = 133;
// bram[3573] = 120;
// bram[3574] = 107;
// bram[3575] = 94;
// bram[3576] = 82;
// bram[3577] = 70;
// bram[3578] = 59;
// bram[3579] = 48;
// bram[3580] = 38;
// bram[3581] = 29;
// bram[3582] = 21;
// bram[3583] = 15;
// bram[3584] = 9;
// bram[3585] = 5;
// bram[3586] = 2;
// bram[3587] = 0;
// bram[3588] = 0;
// bram[3589] = 0;
// bram[3590] = 3;
// bram[3591] = 6;
// bram[3592] = 11;
// bram[3593] = 17;
// bram[3594] = 25;
// bram[3595] = 33;
// bram[3596] = 42;
// bram[3597] = 52;
// bram[3598] = 63;
// bram[3599] = 75;
// bram[3600] = 87;
// bram[3601] = 100;
// bram[3602] = 113;
// bram[3603] = 126;
// bram[3604] = 139;
// bram[3605] = 152;
// bram[3606] = 164;
// bram[3607] = 177;
// bram[3608] = 188;
// bram[3609] = 199;
// bram[3610] = 210;
// bram[3611] = 219;
// bram[3612] = 228;
// bram[3613] = 235;
// bram[3614] = 241;
// bram[3615] = 246;
// bram[3616] = 250;
// bram[3617] = 252;
// bram[3618] = 253;
// bram[3619] = 253;
// bram[3620] = 252;
// bram[3621] = 249;
// bram[3622] = 245;
// bram[3623] = 239;
// bram[3624] = 232;
// bram[3625] = 225;
// bram[3626] = 216;
// bram[3627] = 206;
// bram[3628] = 196;
// bram[3629] = 184;
// bram[3630] = 172;
// bram[3631] = 160;
// bram[3632] = 147;
// bram[3633] = 134;
// bram[3634] = 121;
// bram[3635] = 108;
// bram[3636] = 95;
// bram[3637] = 83;
// bram[3638] = 71;
// bram[3639] = 59;
// bram[3640] = 49;
// bram[3641] = 39;
// bram[3642] = 30;
// bram[3643] = 22;
// bram[3644] = 15;
// bram[3645] = 9;
// bram[3646] = 5;
// bram[3647] = 2;
// bram[3648] = 0;
// bram[3649] = 0;
// bram[3650] = 0;
// bram[3651] = 3;
// bram[3652] = 6;
// bram[3653] = 11;
// bram[3654] = 17;
// bram[3655] = 24;
// bram[3656] = 32;
// bram[3657] = 42;
// bram[3658] = 52;
// bram[3659] = 63;
// bram[3660] = 74;
// bram[3661] = 86;
// bram[3662] = 99;
// bram[3663] = 112;
// bram[3664] = 125;
// bram[3665] = 138;
// bram[3666] = 151;
// bram[3667] = 164;
// bram[3668] = 176;
// bram[3669] = 188;
// bram[3670] = 199;
// bram[3671] = 209;
// bram[3672] = 219;
// bram[3673] = 227;
// bram[3674] = 234;
// bram[3675] = 241;
// bram[3676] = 246;
// bram[3677] = 250;
// bram[3678] = 252;
// bram[3679] = 253;
// bram[3680] = 253;
// bram[3681] = 252;
// bram[3682] = 249;
// bram[3683] = 245;
// bram[3684] = 239;
// bram[3685] = 233;
// bram[3686] = 225;
// bram[3687] = 217;
// bram[3688] = 207;
// bram[3689] = 196;
// bram[3690] = 185;
// bram[3691] = 173;
// bram[3692] = 161;
// bram[3693] = 148;
// bram[3694] = 135;
// bram[3695] = 122;
// bram[3696] = 109;
// bram[3697] = 96;
// bram[3698] = 84;
// bram[3699] = 72;
// bram[3700] = 60;
// bram[3701] = 49;
// bram[3702] = 39;
// bram[3703] = 30;
// bram[3704] = 22;
// bram[3705] = 15;
// bram[3706] = 10;
// bram[3707] = 5;
// bram[3708] = 2;
// bram[3709] = 0;
// bram[3710] = 0;
// bram[3711] = 0;
// bram[3712] = 2;
// bram[3713] = 6;
// bram[3714] = 11;
// bram[3715] = 16;
// bram[3716] = 24;
// bram[3717] = 32;
// bram[3718] = 41;
// bram[3719] = 51;
// bram[3720] = 62;
// bram[3721] = 73;
// bram[3722] = 86;
// bram[3723] = 98;
// bram[3724] = 111;
// bram[3725] = 124;
// bram[3726] = 137;
// bram[3727] = 150;
// bram[3728] = 163;
// bram[3729] = 175;
// bram[3730] = 187;
// bram[3731] = 198;
// bram[3732] = 208;
// bram[3733] = 218;
// bram[3734] = 226;
// bram[3735] = 234;
// bram[3736] = 240;
// bram[3737] = 246;
// bram[3738] = 249;
// bram[3739] = 252;
// bram[3740] = 253;
// bram[3741] = 253;
// bram[3742] = 252;
// bram[3743] = 249;
// bram[3744] = 245;
// bram[3745] = 240;
// bram[3746] = 233;
// bram[3747] = 226;
// bram[3748] = 217;
// bram[3749] = 208;
// bram[3750] = 197;
// bram[3751] = 186;
// bram[3752] = 174;
// bram[3753] = 162;
// bram[3754] = 149;
// bram[3755] = 136;
// bram[3756] = 123;
// bram[3757] = 110;
// bram[3758] = 97;
// bram[3759] = 85;
// bram[3760] = 72;
// bram[3761] = 61;
// bram[3762] = 50;
// bram[3763] = 40;
// bram[3764] = 31;
// bram[3765] = 23;
// bram[3766] = 16;
// bram[3767] = 10;
// bram[3768] = 5;
// bram[3769] = 2;
// bram[3770] = 0;
// bram[3771] = 0;
// bram[3772] = 0;
// bram[3773] = 2;
// bram[3774] = 6;
// bram[3775] = 10;
// bram[3776] = 16;
// bram[3777] = 23;
// bram[3778] = 31;
// bram[3779] = 40;
// bram[3780] = 50;
// bram[3781] = 61;
// bram[3782] = 73;
// bram[3783] = 85;
// bram[3784] = 97;
// bram[3785] = 110;
// bram[3786] = 123;
// bram[3787] = 136;
// bram[3788] = 149;
// bram[3789] = 162;
// bram[3790] = 174;
// bram[3791] = 186;
// bram[3792] = 197;
// bram[3793] = 208;
// bram[3794] = 217;
// bram[3795] = 226;
// bram[3796] = 234;
// bram[3797] = 240;
// bram[3798] = 245;
// bram[3799] = 249;
// bram[3800] = 252;
// bram[3801] = 253;
// bram[3802] = 253;
// bram[3803] = 252;
// bram[3804] = 249;
// bram[3805] = 245;
// bram[3806] = 240;
// bram[3807] = 234;
// bram[3808] = 226;
// bram[3809] = 218;
// bram[3810] = 208;
// bram[3811] = 198;
// bram[3812] = 187;
// bram[3813] = 175;
// bram[3814] = 163;
// bram[3815] = 150;
// bram[3816] = 137;
// bram[3817] = 124;
// bram[3818] = 111;
// bram[3819] = 98;
// bram[3820] = 85;
// bram[3821] = 73;
// bram[3822] = 62;
// bram[3823] = 51;
// bram[3824] = 41;
// bram[3825] = 32;
// bram[3826] = 23;
// bram[3827] = 16;
// bram[3828] = 10;
// bram[3829] = 6;
// bram[3830] = 2;
// bram[3831] = 0;
// bram[3832] = 0;
// bram[3833] = 0;
// bram[3834] = 2;
// bram[3835] = 5;
// bram[3836] = 10;
// bram[3837] = 16;
// bram[3838] = 22;
// bram[3839] = 31;
// bram[3840] = 40;
// bram[3841] = 50;
// bram[3842] = 60;
// bram[3843] = 72;
// bram[3844] = 84;
// bram[3845] = 96;
// bram[3846] = 109;
// bram[3847] = 122;
// bram[3848] = 135;
// bram[3849] = 148;
// bram[3850] = 161;
// bram[3851] = 173;
// bram[3852] = 185;
// bram[3853] = 196;
// bram[3854] = 207;
// bram[3855] = 217;
// bram[3856] = 225;
// bram[3857] = 233;
// bram[3858] = 240;
// bram[3859] = 245;
// bram[3860] = 249;
// bram[3861] = 252;
// bram[3862] = 253;
// bram[3863] = 253;
// bram[3864] = 252;
// bram[3865] = 250;
// bram[3866] = 246;
// bram[3867] = 241;
// bram[3868] = 234;
// bram[3869] = 227;
// bram[3870] = 218;
// bram[3871] = 209;
// bram[3872] = 199;
// bram[3873] = 187;
// bram[3874] = 176;
// bram[3875] = 163;
// bram[3876] = 151;
// bram[3877] = 138;
// bram[3878] = 125;
// bram[3879] = 112;
// bram[3880] = 99;
// bram[3881] = 86;
// bram[3882] = 74;
// bram[3883] = 62;
// bram[3884] = 52;
// bram[3885] = 41;
// bram[3886] = 32;
// bram[3887] = 24;
// bram[3888] = 17;
// bram[3889] = 11;
// bram[3890] = 6;
// bram[3891] = 3;
// bram[3892] = 0;
// bram[3893] = 0;
// bram[3894] = 0;
// bram[3895] = 2;
// bram[3896] = 5;
// bram[3897] = 9;
// bram[3898] = 15;
// bram[3899] = 22;
// bram[3900] = 30;
// bram[3901] = 39;
// bram[3902] = 49;
// bram[3903] = 60;
// bram[3904] = 71;
// bram[3905] = 83;
// bram[3906] = 95;
// bram[3907] = 108;
// bram[3908] = 121;
// bram[3909] = 134;
// bram[3910] = 147;
// bram[3911] = 160;
// bram[3912] = 173;
// bram[3913] = 184;
// bram[3914] = 196;
// bram[3915] = 206;
// bram[3916] = 216;
// bram[3917] = 225;
// bram[3918] = 233;
// bram[3919] = 239;
// bram[3920] = 245;
// bram[3921] = 249;
// bram[3922] = 252;
// bram[3923] = 253;
// bram[3924] = 253;
// bram[3925] = 252;
// bram[3926] = 250;
// bram[3927] = 246;
// bram[3928] = 241;
// bram[3929] = 235;
// bram[3930] = 227;
// bram[3931] = 219;
// bram[3932] = 210;
// bram[3933] = 199;
// bram[3934] = 188;
// bram[3935] = 176;
// bram[3936] = 164;
// bram[3937] = 152;
// bram[3938] = 139;
// bram[3939] = 126;
// bram[3940] = 113;
// bram[3941] = 100;
// bram[3942] = 87;
// bram[3943] = 75;
// bram[3944] = 63;
// bram[3945] = 52;
// bram[3946] = 42;
// bram[3947] = 33;
// bram[3948] = 24;
// bram[3949] = 17;
// bram[3950] = 11;
// bram[3951] = 6;
// bram[3952] = 3;
// bram[3953] = 0;
// bram[3954] = 0;
// bram[3955] = 0;
// bram[3956] = 2;
// bram[3957] = 5;
// bram[3958] = 9;
// bram[3959] = 15;
// bram[3960] = 21;
// bram[3961] = 29;
// bram[3962] = 38;
// bram[3963] = 48;
// bram[3964] = 59;
// bram[3965] = 70;
// bram[3966] = 82;
// bram[3967] = 95;
// bram[3968] = 107;
// bram[3969] = 120;
// bram[3970] = 133;
// bram[3971] = 146;
// bram[3972] = 159;
// bram[3973] = 172;
// bram[3974] = 184;
// bram[3975] = 195;
// bram[3976] = 206;
// bram[3977] = 215;
// bram[3978] = 224;
// bram[3979] = 232;
// bram[3980] = 239;
// bram[3981] = 244;
// bram[3982] = 249;
// bram[3983] = 251;
// bram[3984] = 253;
// bram[3985] = 253;
// bram[3986] = 252;
// bram[3987] = 250;
// bram[3988] = 246;
// bram[3989] = 241;
// bram[3990] = 235;
// bram[3991] = 228;
// bram[3992] = 220;
// bram[3993] = 210;
// bram[3994] = 200;
// bram[3995] = 189;
// bram[3996] = 177;
// bram[3997] = 165;
// bram[3998] = 152;
// bram[3999] = 140;
// bram[4000] = 126;
// bram[4001] = 113;
// bram[4002] = 101;
// bram[4003] = 88;
// bram[4004] = 76;
// bram[4005] = 64;
// bram[4006] = 53;
// bram[4007] = 43;
// bram[4008] = 33;
// bram[4009] = 25;
// bram[4010] = 18;
// bram[4011] = 12;
// bram[4012] = 7;
// bram[4013] = 3;
// bram[4014] = 1;
// bram[4015] = 0;
// bram[4016] = 0;
// bram[4017] = 2;
// bram[4018] = 4;
// bram[4019] = 9;
// bram[4020] = 14;
// bram[4021] = 21;
// bram[4022] = 29;
// bram[4023] = 38;
// bram[4024] = 47;
// bram[4025] = 58;
// bram[4026] = 69;
// bram[4027] = 81;
// bram[4028] = 94;
// bram[4029] = 107;
// bram[4030] = 120;
// bram[4031] = 133;
// bram[4032] = 146;
// bram[4033] = 158;
// bram[4034] = 171;
// bram[4035] = 183;
// bram[4036] = 194;
// bram[4037] = 205;
// bram[4038] = 215;
// bram[4039] = 224;
// bram[4040] = 232;
// bram[4041] = 238;
// bram[4042] = 244;
// bram[4043] = 248;
// bram[4044] = 251;
// bram[4045] = 253;
// bram[4046] = 253;
// bram[4047] = 253;
// bram[4048] = 250;
// bram[4049] = 247;
// bram[4050] = 242;
// bram[4051] = 236;
// bram[4052] = 229;
// bram[4053] = 220;
// bram[4054] = 211;
// bram[4055] = 201;
// bram[4056] = 190;
// bram[4057] = 178;
// bram[4058] = 166;
// bram[4059] = 153;
// bram[4060] = 140;
// bram[4061] = 127;
// bram[4062] = 114;
// bram[4063] = 101;
// bram[4064] = 89;
// bram[4065] = 77;
// bram[4066] = 65;
// bram[4067] = 54;
// bram[4068] = 43;
// bram[4069] = 34;
// bram[4070] = 26;
// bram[4071] = 18;
// bram[4072] = 12;
// bram[4073] = 7;
// bram[4074] = 3;
// bram[4075] = 1;
// bram[4076] = 0;
// bram[4077] = 0;
// bram[4078] = 1;
// bram[4079] = 4;
// bram[4080] = 8;
// bram[4081] = 14;
// bram[4082] = 20;
// bram[4083] = 28;
// bram[4084] = 37;
// bram[4085] = 47;
// bram[4086] = 57;
// bram[4087] = 69;
// bram[4088] = 80;
// bram[4089] = 93;
// bram[4090] = 106;
// bram[4091] = 119;
// bram[4092] = 132;
// bram[4093] = 145;
// bram[4094] = 158;
// bram[4095] = 170;
// bram[4096] = 182;
// bram[4097] = 193;
// bram[4098] = 204;
// bram[4099] = 214;
// bram[4100] = 223;
// bram[4101] = 231;
// bram[4102] = 238;
// bram[4103] = 244;
// bram[4104] = 248;
// bram[4105] = 251;
// bram[4106] = 253;
// bram[4107] = 253;
// bram[4108] = 253;
// bram[4109] = 250;
// bram[4110] = 247;
// bram[4111] = 242;
// bram[4112] = 236;
// bram[4113] = 229;
// bram[4114] = 221;
// bram[4115] = 212;
// bram[4116] = 201;
// bram[4117] = 191;
// bram[4118] = 179;
// bram[4119] = 167;
// bram[4120] = 154;
// bram[4121] = 141;
// bram[4122] = 128;
// bram[4123] = 115;
// bram[4124] = 102;
// bram[4125] = 90;
// bram[4126] = 77;
// bram[4127] = 66;
// bram[4128] = 54;
// bram[4129] = 44;
// bram[4130] = 35;
// bram[4131] = 26;
// bram[4132] = 19;
// bram[4133] = 12;
// bram[4134] = 7;
// bram[4135] = 3;
// bram[4136] = 1;
// bram[4137] = 0;
// bram[4138] = 0;
// bram[4139] = 1;
// bram[4140] = 4;
// bram[4141] = 8;
// bram[4142] = 13;
// bram[4143] = 20;
// bram[4144] = 28;
// bram[4145] = 36;
// bram[4146] = 46;
// bram[4147] = 57;
// bram[4148] = 68;
// bram[4149] = 80;
// bram[4150] = 92;
// bram[4151] = 105;
// bram[4152] = 118;
// bram[4153] = 131;
// bram[4154] = 144;
// bram[4155] = 157;
// bram[4156] = 169;
// bram[4157] = 181;
// bram[4158] = 193;
// bram[4159] = 203;
// bram[4160] = 213;
// bram[4161] = 222;
// bram[4162] = 231;
// bram[4163] = 237;
// bram[4164] = 243;
// bram[4165] = 248;
// bram[4166] = 251;
// bram[4167] = 253;
// bram[4168] = 253;
// bram[4169] = 253;
// bram[4170] = 251;
// bram[4171] = 247;
// bram[4172] = 243;
// bram[4173] = 237;
// bram[4174] = 230;
// bram[4175] = 221;
// bram[4176] = 212;
// bram[4177] = 202;
// bram[4178] = 191;
// bram[4179] = 180;
// bram[4180] = 168;
// bram[4181] = 155;
// bram[4182] = 142;
// bram[4183] = 129;
// bram[4184] = 116;
// bram[4185] = 103;
// bram[4186] = 90;
// bram[4187] = 78;
// bram[4188] = 66;
// bram[4189] = 55;
// bram[4190] = 45;
// bram[4191] = 35;
// bram[4192] = 27;
// bram[4193] = 19;
// bram[4194] = 13;
// bram[4195] = 8;
// bram[4196] = 4;
// bram[4197] = 1;
// bram[4198] = 0;
// bram[4199] = 0;
// bram[4200] = 1;
// bram[4201] = 4;
// bram[4202] = 8;
// bram[4203] = 13;
// bram[4204] = 19;
// bram[4205] = 27;
// bram[4206] = 36;
// bram[4207] = 45;
// bram[4208] = 56;
// bram[4209] = 67;
// bram[4210] = 79;
// bram[4211] = 91;
// bram[4212] = 104;
// bram[4213] = 117;
// bram[4214] = 130;
// bram[4215] = 143;
// bram[4216] = 156;
// bram[4217] = 168;
// bram[4218] = 180;
// bram[4219] = 192;
// bram[4220] = 203;
// bram[4221] = 213;
// bram[4222] = 222;
// bram[4223] = 230;
// bram[4224] = 237;
// bram[4225] = 243;
// bram[4226] = 247;
// bram[4227] = 251;
// bram[4228] = 253;
// bram[4229] = 253;
// bram[4230] = 253;
// bram[4231] = 251;
// bram[4232] = 248;
// bram[4233] = 243;
// bram[4234] = 237;
// bram[4235] = 230;
// bram[4236] = 222;
// bram[4237] = 213;
// bram[4238] = 203;
// bram[4239] = 192;
// bram[4240] = 181;
// bram[4241] = 168;
// bram[4242] = 156;
// bram[4243] = 143;
// bram[4244] = 130;
// bram[4245] = 117;
// bram[4246] = 104;
// bram[4247] = 91;
// bram[4248] = 79;
// bram[4249] = 67;
// bram[4250] = 56;
// bram[4251] = 45;
// bram[4252] = 36;
// bram[4253] = 27;
// bram[4254] = 20;
// bram[4255] = 13;
// bram[4256] = 8;
// bram[4257] = 4;
// bram[4258] = 1;
// bram[4259] = 0;
// bram[4260] = 0;
// bram[4261] = 1;
// bram[4262] = 4;
// bram[4263] = 7;
// bram[4264] = 13;
// bram[4265] = 19;
// bram[4266] = 27;
// bram[4267] = 35;
// bram[4268] = 45;
// bram[4269] = 55;
// bram[4270] = 66;
// bram[4271] = 78;
// bram[4272] = 90;
// bram[4273] = 103;
// bram[4274] = 116;
// bram[4275] = 129;
// bram[4276] = 142;
// bram[4277] = 155;
// bram[4278] = 167;
// bram[4279] = 180;
// bram[4280] = 191;
// bram[4281] = 202;
// bram[4282] = 212;
// bram[4283] = 221;
// bram[4284] = 229;
// bram[4285] = 237;
// bram[4286] = 242;
// bram[4287] = 247;
// bram[4288] = 251;
// bram[4289] = 253;
// bram[4290] = 253;
// bram[4291] = 253;
// bram[4292] = 251;
// bram[4293] = 248;
// bram[4294] = 243;
// bram[4295] = 238;
// bram[4296] = 231;
// bram[4297] = 223;
// bram[4298] = 214;
// bram[4299] = 204;
// bram[4300] = 193;
// bram[4301] = 181;
// bram[4302] = 169;
// bram[4303] = 157;
// bram[4304] = 144;
// bram[4305] = 131;
// bram[4306] = 118;
// bram[4307] = 105;
// bram[4308] = 92;
// bram[4309] = 80;
// bram[4310] = 68;
// bram[4311] = 57;
// bram[4312] = 46;
// bram[4313] = 36;
// bram[4314] = 28;
// bram[4315] = 20;
// bram[4316] = 14;
// bram[4317] = 8;
// bram[4318] = 4;
// bram[4319] = 1;
// bram[4320] = 0;
// bram[4321] = 0;
// bram[4322] = 1;
// bram[4323] = 3;
// bram[4324] = 7;
// bram[4325] = 12;
// bram[4326] = 19;
// bram[4327] = 26;
// bram[4328] = 34;
// bram[4329] = 44;
// bram[4330] = 54;
// bram[4331] = 65;
// bram[4332] = 77;
// bram[4333] = 89;
// bram[4334] = 102;
// bram[4335] = 115;
// bram[4336] = 128;
// bram[4337] = 141;
// bram[4338] = 154;
// bram[4339] = 167;
// bram[4340] = 179;
// bram[4341] = 190;
// bram[4342] = 201;
// bram[4343] = 211;
// bram[4344] = 221;
// bram[4345] = 229;
// bram[4346] = 236;
// bram[4347] = 242;
// bram[4348] = 247;
// bram[4349] = 250;
// bram[4350] = 253;
// bram[4351] = 253;
// bram[4352] = 253;
// bram[4353] = 251;
// bram[4354] = 248;
// bram[4355] = 244;
// bram[4356] = 238;
// bram[4357] = 231;
// bram[4358] = 223;
// bram[4359] = 214;
// bram[4360] = 204;
// bram[4361] = 194;
// bram[4362] = 182;
// bram[4363] = 170;
// bram[4364] = 158;
// bram[4365] = 145;
// bram[4366] = 132;
// bram[4367] = 119;
// bram[4368] = 106;
// bram[4369] = 93;
// bram[4370] = 81;
// bram[4371] = 69;
// bram[4372] = 57;
// bram[4373] = 47;
// bram[4374] = 37;
// bram[4375] = 28;
// bram[4376] = 21;
// bram[4377] = 14;
// bram[4378] = 8;
// bram[4379] = 4;
// bram[4380] = 1;
// bram[4381] = 0;
// bram[4382] = 0;
// bram[4383] = 1;
// bram[4384] = 3;
// bram[4385] = 7;
// bram[4386] = 12;
// bram[4387] = 18;
// bram[4388] = 25;
// bram[4389] = 34;
// bram[4390] = 43;
// bram[4391] = 54;
// bram[4392] = 65;
// bram[4393] = 76;
// bram[4394] = 89;
// bram[4395] = 101;
// bram[4396] = 114;
// bram[4397] = 127;
// bram[4398] = 140;
// bram[4399] = 153;
// bram[4400] = 166;
// bram[4401] = 178;
// bram[4402] = 190;
// bram[4403] = 201;
// bram[4404] = 211;
// bram[4405] = 220;
// bram[4406] = 228;
// bram[4407] = 236;
// bram[4408] = 242;
// bram[4409] = 247;
// bram[4410] = 250;
// bram[4411] = 253;
// bram[4412] = 253;
// bram[4413] = 253;
// bram[4414] = 251;
// bram[4415] = 248;
// bram[4416] = 244;
// bram[4417] = 238;
// bram[4418] = 232;
// bram[4419] = 224;
// bram[4420] = 215;
// bram[4421] = 205;
// bram[4422] = 194;
// bram[4423] = 183;
// bram[4424] = 171;
// bram[4425] = 159;
// bram[4426] = 146;
// bram[4427] = 133;
// bram[4428] = 120;
// bram[4429] = 107;
// bram[4430] = 94;
// bram[4431] = 82;
// bram[4432] = 70;
// bram[4433] = 58;
// bram[4434] = 48;
// bram[4435] = 38;
// bram[4436] = 29;
// bram[4437] = 21;
// bram[4438] = 14;
// bram[4439] = 9;
// bram[4440] = 5;
// bram[4441] = 2;
// bram[4442] = 0;
// bram[4443] = 0;
// bram[4444] = 1;
// bram[4445] = 3;
// bram[4446] = 7;
// bram[4447] = 11;
// bram[4448] = 18;
// bram[4449] = 25;
// bram[4450] = 33;
// bram[4451] = 43;
// bram[4452] = 53;
// bram[4453] = 64;
// bram[4454] = 76;
// bram[4455] = 88;
// bram[4456] = 100;
// bram[4457] = 113;
// bram[4458] = 126;
// bram[4459] = 139;
// bram[4460] = 152;
// bram[4461] = 165;
// bram[4462] = 177;
// bram[4463] = 189;
// bram[4464] = 200;
// bram[4465] = 210;
// bram[4466] = 219;
// bram[4467] = 228;
// bram[4468] = 235;
// bram[4469] = 241;
// bram[4470] = 246;
// bram[4471] = 250;
// bram[4472] = 252;
// bram[4473] = 253;
// bram[4474] = 253;
// bram[4475] = 252;
// bram[4476] = 249;
// bram[4477] = 244;
// bram[4478] = 239;
// bram[4479] = 232;
// bram[4480] = 224;
// bram[4481] = 216;
// bram[4482] = 206;
// bram[4483] = 195;
// bram[4484] = 184;
// bram[4485] = 172;
// bram[4486] = 159;
// bram[4487] = 147;
// bram[4488] = 134;
// bram[4489] = 121;
// bram[4490] = 108;
// bram[4491] = 95;
// bram[4492] = 82;
// bram[4493] = 70;
// bram[4494] = 59;
// bram[4495] = 48;
// bram[4496] = 38;
// bram[4497] = 29;
// bram[4498] = 22;
// bram[4499] = 15;
// bram[4500] = 9;
// bram[4501] = 5;
// bram[4502] = 2;
// bram[4503] = 0;
// bram[4504] = 0;
// bram[4505] = 0;
// bram[4506] = 3;
// bram[4507] = 6;
// bram[4508] = 11;
// bram[4509] = 17;
// bram[4510] = 24;
// bram[4511] = 33;
// bram[4512] = 42;
// bram[4513] = 52;
// bram[4514] = 63;
// bram[4515] = 75;
// bram[4516] = 87;
// bram[4517] = 99;
// bram[4518] = 112;
// bram[4519] = 125;
// bram[4520] = 138;
// bram[4521] = 151;
// bram[4522] = 164;
// bram[4523] = 176;
// bram[4524] = 188;
// bram[4525] = 199;
// bram[4526] = 209;
// bram[4527] = 219;
// bram[4528] = 227;
// bram[4529] = 235;
// bram[4530] = 241;
// bram[4531] = 246;
// bram[4532] = 250;
// bram[4533] = 252;
// bram[4534] = 253;
// bram[4535] = 253;
// bram[4536] = 252;
// bram[4537] = 249;
// bram[4538] = 245;
// bram[4539] = 239;
// bram[4540] = 233;
// bram[4541] = 225;
// bram[4542] = 216;
// bram[4543] = 206;
// bram[4544] = 196;
// bram[4545] = 185;
// bram[4546] = 173;
// bram[4547] = 160;
// bram[4548] = 148;
// bram[4549] = 135;
// bram[4550] = 122;
// bram[4551] = 109;
// bram[4552] = 96;
// bram[4553] = 83;
// bram[4554] = 71;
// bram[4555] = 60;
// bram[4556] = 49;
// bram[4557] = 39;
// bram[4558] = 30;
// bram[4559] = 22;
// bram[4560] = 15;
// bram[4561] = 10;
// bram[4562] = 5;
// bram[4563] = 2;
// bram[4564] = 0;
// bram[4565] = 0;
// bram[4566] = 0;
// bram[4567] = 2;
// bram[4568] = 6;
// bram[4569] = 11;
// bram[4570] = 17;
// bram[4571] = 24;
// bram[4572] = 32;
// bram[4573] = 41;
// bram[4574] = 51;
// bram[4575] = 62;
// bram[4576] = 74;
// bram[4577] = 86;
// bram[4578] = 99;
// bram[4579] = 111;
// bram[4580] = 125;
// bram[4581] = 138;
// bram[4582] = 150;
// bram[4583] = 163;
// bram[4584] = 175;
// bram[4585] = 187;
// bram[4586] = 198;
// bram[4587] = 209;
// bram[4588] = 218;
// bram[4589] = 227;
// bram[4590] = 234;
// bram[4591] = 241;
// bram[4592] = 246;
// bram[4593] = 250;
// bram[4594] = 252;
// bram[4595] = 253;
// bram[4596] = 253;
// bram[4597] = 252;
// bram[4598] = 249;
// bram[4599] = 245;
// bram[4600] = 240;
// bram[4601] = 233;
// bram[4602] = 225;
// bram[4603] = 217;
// bram[4604] = 207;
// bram[4605] = 197;
// bram[4606] = 185;
// bram[4607] = 174;
// bram[4608] = 161;
// bram[4609] = 148;
// bram[4610] = 135;
// bram[4611] = 122;
// bram[4612] = 109;
// bram[4613] = 97;
// bram[4614] = 84;
// bram[4615] = 72;
// bram[4616] = 60;
// bram[4617] = 50;
// bram[4618] = 40;
// bram[4619] = 31;
// bram[4620] = 23;
// bram[4621] = 16;
// bram[4622] = 10;
// bram[4623] = 5;
// bram[4624] = 2;
// bram[4625] = 0;
// bram[4626] = 0;
// bram[4627] = 0;
// bram[4628] = 2;
// bram[4629] = 6;
// bram[4630] = 10;
// bram[4631] = 16;
// bram[4632] = 23;
// bram[4633] = 31;
// bram[4634] = 41;
// bram[4635] = 51;
// bram[4636] = 62;
// bram[4637] = 73;
// bram[4638] = 85;
// bram[4639] = 98;
// bram[4640] = 111;
// bram[4641] = 124;
// bram[4642] = 137;
// bram[4643] = 150;
// bram[4644] = 162;
// bram[4645] = 175;
// bram[4646] = 186;
// bram[4647] = 198;
// bram[4648] = 208;
// bram[4649] = 218;
// bram[4650] = 226;
// bram[4651] = 234;
// bram[4652] = 240;
// bram[4653] = 245;
// bram[4654] = 249;
// bram[4655] = 252;
// bram[4656] = 253;
// bram[4657] = 253;
// bram[4658] = 252;
// bram[4659] = 249;
// bram[4660] = 245;
// bram[4661] = 240;
// bram[4662] = 234;
// bram[4663] = 226;
// bram[4664] = 217;
// bram[4665] = 208;
// bram[4666] = 197;
// bram[4667] = 186;
// bram[4668] = 174;
// bram[4669] = 162;
// bram[4670] = 149;
// bram[4671] = 136;
// bram[4672] = 123;
// bram[4673] = 110;
// bram[4674] = 97;
// bram[4675] = 85;
// bram[4676] = 73;
// bram[4677] = 61;
// bram[4678] = 50;
// bram[4679] = 40;
// bram[4680] = 31;
// bram[4681] = 23;
// bram[4682] = 16;
// bram[4683] = 10;
// bram[4684] = 6;
// bram[4685] = 2;
// bram[4686] = 0;
// bram[4687] = 0;
// bram[4688] = 0;
// bram[4689] = 2;
// bram[4690] = 5;
// bram[4691] = 10;
// bram[4692] = 16;
// bram[4693] = 23;
// bram[4694] = 31;
// bram[4695] = 40;
// bram[4696] = 50;
// bram[4697] = 61;
// bram[4698] = 72;
// bram[4699] = 84;
// bram[4700] = 97;
// bram[4701] = 110;
// bram[4702] = 123;
// bram[4703] = 136;
// bram[4704] = 149;
// bram[4705] = 161;
// bram[4706] = 174;
// bram[4707] = 186;
// bram[4708] = 197;
// bram[4709] = 207;
// bram[4710] = 217;
// bram[4711] = 226;
// bram[4712] = 233;
// bram[4713] = 240;
// bram[4714] = 245;
// bram[4715] = 249;
// bram[4716] = 252;
// bram[4717] = 253;
// bram[4718] = 253;
// bram[4719] = 252;
// bram[4720] = 250;
// bram[4721] = 246;
// bram[4722] = 240;
// bram[4723] = 234;
// bram[4724] = 227;
// bram[4725] = 218;
// bram[4726] = 209;
// bram[4727] = 198;
// bram[4728] = 187;
// bram[4729] = 175;
// bram[4730] = 163;
// bram[4731] = 150;
// bram[4732] = 137;
// bram[4733] = 124;
// bram[4734] = 111;
// bram[4735] = 98;
// bram[4736] = 86;
// bram[4737] = 74;
// bram[4738] = 62;
// bram[4739] = 51;
// bram[4740] = 41;
// bram[4741] = 32;
// bram[4742] = 24;
// bram[4743] = 17;
// bram[4744] = 11;
// bram[4745] = 6;
// bram[4746] = 2;
// bram[4747] = 0;
// bram[4748] = 0;
// bram[4749] = 0;
// bram[4750] = 2;
// bram[4751] = 5;
// bram[4752] = 10;
// bram[4753] = 15;
// bram[4754] = 22;
// bram[4755] = 30;
// bram[4756] = 39;
// bram[4757] = 49;
// bram[4758] = 60;
// bram[4759] = 71;
// bram[4760] = 83;
// bram[4761] = 96;
// bram[4762] = 109;
// bram[4763] = 122;
// bram[4764] = 135;
// bram[4765] = 148;
// bram[4766] = 161;
// bram[4767] = 173;
// bram[4768] = 185;
// bram[4769] = 196;
// bram[4770] = 207;
// bram[4771] = 216;
// bram[4772] = 225;
// bram[4773] = 233;
// bram[4774] = 239;
// bram[4775] = 245;
// bram[4776] = 249;
// bram[4777] = 252;
// bram[4778] = 253;
// bram[4779] = 253;
// bram[4780] = 252;
// bram[4781] = 250;
// bram[4782] = 246;
// bram[4783] = 241;
// bram[4784] = 235;
// bram[4785] = 227;
// bram[4786] = 219;
// bram[4787] = 209;
// bram[4788] = 199;
// bram[4789] = 188;
// bram[4790] = 176;
// bram[4791] = 164;
// bram[4792] = 151;
// bram[4793] = 138;
// bram[4794] = 125;
// bram[4795] = 112;
// bram[4796] = 99;
// bram[4797] = 87;
// bram[4798] = 74;
// bram[4799] = 63;
// bram[4800] = 52;
// bram[4801] = 42;
// bram[4802] = 32;
// bram[4803] = 24;
// bram[4804] = 17;
// bram[4805] = 11;
// bram[4806] = 6;
// bram[4807] = 3;
// bram[4808] = 0;
// bram[4809] = 0;
// bram[4810] = 0;
// bram[4811] = 2;
// bram[4812] = 5;
// bram[4813] = 9;
// bram[4814] = 15;
// bram[4815] = 22;
// bram[4816] = 30;
// bram[4817] = 39;
// bram[4818] = 49;
// bram[4819] = 59;
// bram[4820] = 71;
// bram[4821] = 83;
// bram[4822] = 95;
// bram[4823] = 108;
// bram[4824] = 121;
// bram[4825] = 134;
// bram[4826] = 147;
// bram[4827] = 160;
// bram[4828] = 172;
// bram[4829] = 184;
// bram[4830] = 195;
// bram[4831] = 206;
// bram[4832] = 216;
// bram[4833] = 225;
// bram[4834] = 232;
// bram[4835] = 239;
// bram[4836] = 244;
// bram[4837] = 249;
// bram[4838] = 252;
// bram[4839] = 253;
// bram[4840] = 253;
// bram[4841] = 252;
// bram[4842] = 250;
// bram[4843] = 246;
// bram[4844] = 241;
// bram[4845] = 235;
// bram[4846] = 228;
// bram[4847] = 219;
// bram[4848] = 210;
// bram[4849] = 200;
// bram[4850] = 189;
// bram[4851] = 177;
// bram[4852] = 165;
// bram[4853] = 152;
// bram[4854] = 139;
// bram[4855] = 126;
// bram[4856] = 113;
// bram[4857] = 100;
// bram[4858] = 87;
// bram[4859] = 75;
// bram[4860] = 64;
// bram[4861] = 53;
// bram[4862] = 42;
// bram[4863] = 33;
// bram[4864] = 25;
// bram[4865] = 17;
// bram[4866] = 11;
// bram[4867] = 6;
// bram[4868] = 3;
// bram[4869] = 1;
// bram[4870] = 0;
// bram[4871] = 0;
// bram[4872] = 2;
// bram[4873] = 5;
// bram[4874] = 9;
// bram[4875] = 14;
// bram[4876] = 21;
// bram[4877] = 29;
// bram[4878] = 38;
// bram[4879] = 48;
// bram[4880] = 58;
// bram[4881] = 70;
// bram[4882] = 82;
// bram[4883] = 94;
// bram[4884] = 107;
// bram[4885] = 120;
// bram[4886] = 133;
// bram[4887] = 146;
// bram[4888] = 159;
// bram[4889] = 171;
// bram[4890] = 183;
// bram[4891] = 195;
// bram[4892] = 205;
// bram[4893] = 215;
// bram[4894] = 224;
// bram[4895] = 232;
// bram[4896] = 239;
// bram[4897] = 244;
// bram[4898] = 248;
// bram[4899] = 251;
// bram[4900] = 253;
// bram[4901] = 253;
// bram[4902] = 252;
// bram[4903] = 250;
// bram[4904] = 247;
// bram[4905] = 242;
// bram[4906] = 236;
// bram[4907] = 228;
// bram[4908] = 220;
// bram[4909] = 211;
// bram[4910] = 200;
// bram[4911] = 189;
// bram[4912] = 178;
// bram[4913] = 165;
// bram[4914] = 153;
// bram[4915] = 140;
// bram[4916] = 127;
// bram[4917] = 114;
// bram[4918] = 101;
// bram[4919] = 88;
// bram[4920] = 76;
// bram[4921] = 64;
// bram[4922] = 53;
// bram[4923] = 43;
// bram[4924] = 34;
// bram[4925] = 25;
// bram[4926] = 18;
// bram[4927] = 12;
// bram[4928] = 7;
// bram[4929] = 3;
// bram[4930] = 1;
// bram[4931] = 0;
// bram[4932] = 0;
// bram[4933] = 1;
// bram[4934] = 4;
// bram[4935] = 9;
// bram[4936] = 14;
// bram[4937] = 21;
// bram[4938] = 29;
// bram[4939] = 37;
// bram[4940] = 47;
// bram[4941] = 58;
// bram[4942] = 69;
// bram[4943] = 81;
// bram[4944] = 93;
// bram[4945] = 106;
// bram[4946] = 119;
// bram[4947] = 132;
// bram[4948] = 145;
// bram[4949] = 158;
// bram[4950] = 170;
// bram[4951] = 182;
// bram[4952] = 194;
// bram[4953] = 205;
// bram[4954] = 214;
// bram[4955] = 223;
// bram[4956] = 231;
// bram[4957] = 238;
// bram[4958] = 244;
// bram[4959] = 248;
// bram[4960] = 251;
// bram[4961] = 253;
// bram[4962] = 253;
// bram[4963] = 253;
// bram[4964] = 250;
// bram[4965] = 247;
// bram[4966] = 242;
// bram[4967] = 236;
// bram[4968] = 229;
// bram[4969] = 221;
// bram[4970] = 211;
// bram[4971] = 201;
// bram[4972] = 190;
// bram[4973] = 178;
// bram[4974] = 166;
// bram[4975] = 154;
// bram[4976] = 141;
// bram[4977] = 128;
// bram[4978] = 115;
// bram[4979] = 102;
// bram[4980] = 89;
// bram[4981] = 77;
// bram[4982] = 65;
// bram[4983] = 54;
// bram[4984] = 44;
// bram[4985] = 34;
// bram[4986] = 26;
// bram[4987] = 18;
// bram[4988] = 12;
// bram[4989] = 7;
// bram[4990] = 3;
// bram[4991] = 1;
// bram[4992] = 0;
// bram[4993] = 0;
// bram[4994] = 1;
// bram[4995] = 4;
// bram[4996] = 8;
// bram[4997] = 14;
// bram[4998] = 20;
// bram[4999] = 28;
// bram[5000] = 37;
// bram[5001] = 46;
// bram[5002] = 57;
// bram[5003] = 68;
// bram[5004] = 80;
// bram[5005] = 93;
// bram[5006] = 105;
// bram[5007] = 118;
// bram[5008] = 131;
// bram[5009] = 144;
// bram[5010] = 157;
// bram[5011] = 170;
// bram[5012] = 182;
// bram[5013] = 193;
// bram[5014] = 204;
// bram[5015] = 214;
// bram[5016] = 223;
// bram[5017] = 231;
// bram[5018] = 238;
// bram[5019] = 243;
// bram[5020] = 248;
// bram[5021] = 251;
// bram[5022] = 253;
// bram[5023] = 253;
// bram[5024] = 253;
// bram[5025] = 251;
// bram[5026] = 247;
// bram[5027] = 242;
// bram[5028] = 236;
// bram[5029] = 229;
// bram[5030] = 221;
// bram[5031] = 212;
// bram[5032] = 202;
// bram[5033] = 191;
// bram[5034] = 179;
// bram[5035] = 167;
// bram[5036] = 155;
// bram[5037] = 142;
// bram[5038] = 129;
// bram[5039] = 116;
// bram[5040] = 103;
// bram[5041] = 90;
// bram[5042] = 78;
// bram[5043] = 66;
// bram[5044] = 55;
// bram[5045] = 44;
// bram[5046] = 35;
// bram[5047] = 26;
// bram[5048] = 19;
// bram[5049] = 12;
// bram[5050] = 7;
// bram[5051] = 3;
// bram[5052] = 1;
// bram[5053] = 0;
// bram[5054] = 0;
// bram[5055] = 1;
// bram[5056] = 4;
// bram[5057] = 8;
// bram[5058] = 13;
// bram[5059] = 20;
// bram[5060] = 27;
// bram[5061] = 36;
// bram[5062] = 46;
// bram[5063] = 56;
// bram[5064] = 67;
// bram[5065] = 79;
// bram[5066] = 92;
// bram[5067] = 104;
// bram[5068] = 117;
// bram[5069] = 130;
// bram[5070] = 143;
// bram[5071] = 156;
// bram[5072] = 169;
// bram[5073] = 181;
// bram[5074] = 192;
// bram[5075] = 203;
// bram[5076] = 213;
// bram[5077] = 222;
// bram[5078] = 230;
// bram[5079] = 237;
// bram[5080] = 243;
// bram[5081] = 248;
// bram[5082] = 251;
// bram[5083] = 253;
// bram[5084] = 253;
// bram[5085] = 253;
// bram[5086] = 251;
// bram[5087] = 247;
// bram[5088] = 243;
// bram[5089] = 237;
// bram[5090] = 230;
// bram[5091] = 222;
// bram[5092] = 213;
// bram[5093] = 203;
// bram[5094] = 192;
// bram[5095] = 180;
// bram[5096] = 168;
// bram[5097] = 155;
// bram[5098] = 143;
// bram[5099] = 130;
// bram[5100] = 117;
// bram[5101] = 104;
// bram[5102] = 91;
// bram[5103] = 79;
// bram[5104] = 67;
// bram[5105] = 56;
// bram[5106] = 45;
// bram[5107] = 36;
// bram[5108] = 27;
// bram[5109] = 19;
// bram[5110] = 13;
// bram[5111] = 8;
// bram[5112] = 4;
// bram[5113] = 1;
// bram[5114] = 0;
// bram[5115] = 0;
// bram[5116] = 1;
// bram[5117] = 4;
// bram[5118] = 8;
// bram[5119] = 13;
// bram[5120] = 19;
// bram[5121] = 27;
// bram[5122] = 35;
// bram[5123] = 45;
// bram[5124] = 55;
// bram[5125] = 67;
// bram[5126] = 78;
// bram[5127] = 91;
// bram[5128] = 103;
// bram[5129] = 116;
// bram[5130] = 129;
// bram[5131] = 143;
// bram[5132] = 155;
// bram[5133] = 168;
// bram[5134] = 180;
// bram[5135] = 192;
// bram[5136] = 202;
// bram[5137] = 212;
// bram[5138] = 222;
// bram[5139] = 230;
// bram[5140] = 237;
// bram[5141] = 243;
// bram[5142] = 247;
// bram[5143] = 251;
// bram[5144] = 253;
// bram[5145] = 253;
// bram[5146] = 253;
// bram[5147] = 251;
// bram[5148] = 248;
// bram[5149] = 243;
// bram[5150] = 237;
// bram[5151] = 230;
// bram[5152] = 222;
// bram[5153] = 213;
// bram[5154] = 203;
// bram[5155] = 192;
// bram[5156] = 181;
// bram[5157] = 169;
// bram[5158] = 156;
// bram[5159] = 144;
// bram[5160] = 130;
// bram[5161] = 117;
// bram[5162] = 104;
// bram[5163] = 92;
// bram[5164] = 79;
// bram[5165] = 68;
// bram[5166] = 56;
// bram[5167] = 46;
// bram[5168] = 36;
// bram[5169] = 27;
// bram[5170] = 20;
// bram[5171] = 13;
// bram[5172] = 8;
// bram[5173] = 4;
// bram[5174] = 1;
// bram[5175] = 0;
// bram[5176] = 0;
// bram[5177] = 1;
// bram[5178] = 3;
// bram[5179] = 7;
// bram[5180] = 12;
// bram[5181] = 19;
// bram[5182] = 26;
// bram[5183] = 35;
// bram[5184] = 44;
// bram[5185] = 55;
// bram[5186] = 66;
// bram[5187] = 78;
// bram[5188] = 90;
// bram[5189] = 103;
// bram[5190] = 116;
// bram[5191] = 129;
// bram[5192] = 142;
// bram[5193] = 154;
// bram[5194] = 167;
// bram[5195] = 179;
// bram[5196] = 191;
// bram[5197] = 202;
// bram[5198] = 212;
// bram[5199] = 221;
// bram[5200] = 229;
// bram[5201] = 236;
// bram[5202] = 242;
// bram[5203] = 247;
// bram[5204] = 251;
// bram[5205] = 253;
// bram[5206] = 253;
// bram[5207] = 253;
// bram[5208] = 251;
// bram[5209] = 248;
// bram[5210] = 243;
// bram[5211] = 238;
// bram[5212] = 231;
// bram[5213] = 223;
// bram[5214] = 214;
// bram[5215] = 204;
// bram[5216] = 193;
// bram[5217] = 182;
// bram[5218] = 170;
// bram[5219] = 157;
// bram[5220] = 144;
// bram[5221] = 131;
// bram[5222] = 118;
// bram[5223] = 105;
// bram[5224] = 93;
// bram[5225] = 80;
// bram[5226] = 68;
// bram[5227] = 57;
// bram[5228] = 46;
// bram[5229] = 37;
// bram[5230] = 28;
// bram[5231] = 20;
// bram[5232] = 14;
// bram[5233] = 8;
// bram[5234] = 4;
// bram[5235] = 1;
// bram[5236] = 0;
// bram[5237] = 0;
// bram[5238] = 1;
// bram[5239] = 3;
// bram[5240] = 7;
// bram[5241] = 12;
// bram[5242] = 18;
// bram[5243] = 26;
// bram[5244] = 34;
// bram[5245] = 44;
// bram[5246] = 54;
// bram[5247] = 65;
// bram[5248] = 77;
// bram[5249] = 89;
// bram[5250] = 102;
// bram[5251] = 115;
// bram[5252] = 128;
// bram[5253] = 141;
// bram[5254] = 154;
// bram[5255] = 166;
// bram[5256] = 178;
// bram[5257] = 190;
// bram[5258] = 201;
// bram[5259] = 211;
// bram[5260] = 220;
// bram[5261] = 229;
// bram[5262] = 236;
// bram[5263] = 242;
// bram[5264] = 247;
// bram[5265] = 250;
// bram[5266] = 253;
// bram[5267] = 253;
// bram[5268] = 253;
// bram[5269] = 251;
// bram[5270] = 248;
// bram[5271] = 244;
// bram[5272] = 238;
// bram[5273] = 231;
// bram[5274] = 223;
// bram[5275] = 215;
// bram[5276] = 205;
// bram[5277] = 194;
// bram[5278] = 183;
// bram[5279] = 171;
// bram[5280] = 158;
// bram[5281] = 145;
// bram[5282] = 132;
// bram[5283] = 119;
// bram[5284] = 106;
// bram[5285] = 93;
// bram[5286] = 81;
// bram[5287] = 69;
// bram[5288] = 58;
// bram[5289] = 47;
// bram[5290] = 37;
// bram[5291] = 29;
// bram[5292] = 21;
// bram[5293] = 14;
// bram[5294] = 9;
// bram[5295] = 4;
// bram[5296] = 1;
// bram[5297] = 0;
// bram[5298] = 0;
// bram[5299] = 1;
// bram[5300] = 3;
// bram[5301] = 7;
// bram[5302] = 12;
// bram[5303] = 18;
// bram[5304] = 25;
// bram[5305] = 34;
// bram[5306] = 43;
// bram[5307] = 53;
// bram[5308] = 64;
// bram[5309] = 76;
// bram[5310] = 88;
// bram[5311] = 101;
// bram[5312] = 114;
// bram[5313] = 127;
// bram[5314] = 140;
// bram[5315] = 153;
// bram[5316] = 165;
// bram[5317] = 178;
// bram[5318] = 189;
// bram[5319] = 200;
// bram[5320] = 210;
// bram[5321] = 220;
// bram[5322] = 228;
// bram[5323] = 235;
// bram[5324] = 242;
// bram[5325] = 246;
// bram[5326] = 250;
// bram[5327] = 252;
// bram[5328] = 253;
// bram[5329] = 253;
// bram[5330] = 251;
// bram[5331] = 248;
// bram[5332] = 244;
// bram[5333] = 239;
// bram[5334] = 232;
// bram[5335] = 224;
// bram[5336] = 215;
// bram[5337] = 205;
// bram[5338] = 195;
// bram[5339] = 183;
// bram[5340] = 171;
// bram[5341] = 159;
// bram[5342] = 146;
// bram[5343] = 133;
// bram[5344] = 120;
// bram[5345] = 107;
// bram[5346] = 94;
// bram[5347] = 82;
// bram[5348] = 70;
// bram[5349] = 59;
// bram[5350] = 48;
// bram[5351] = 38;
// bram[5352] = 29;
// bram[5353] = 21;
// bram[5354] = 15;
// bram[5355] = 9;
// bram[5356] = 5;
// bram[5357] = 2;
// bram[5358] = 0;
// bram[5359] = 0;
// bram[5360] = 1;
// bram[5361] = 3;
// bram[5362] = 6;
// bram[5363] = 11;
// bram[5364] = 17;
// bram[5365] = 25;
// bram[5366] = 33;
// bram[5367] = 42;
// bram[5368] = 52;
// bram[5369] = 63;
// bram[5370] = 75;
// bram[5371] = 87;
// bram[5372] = 100;
// bram[5373] = 113;
// bram[5374] = 126;
// bram[5375] = 139;
// bram[5376] = 152;
// bram[5377] = 165;
// bram[5378] = 177;
// bram[5379] = 188;
// bram[5380] = 200;
// bram[5381] = 210;
// bram[5382] = 219;
// bram[5383] = 228;
// bram[5384] = 235;
// bram[5385] = 241;
// bram[5386] = 246;
// bram[5387] = 250;
// bram[5388] = 252;
// bram[5389] = 253;
// bram[5390] = 253;
// bram[5391] = 252;
// bram[5392] = 249;
// bram[5393] = 244;
// bram[5394] = 239;
// bram[5395] = 232;
// bram[5396] = 225;
// bram[5397] = 216;
// bram[5398] = 206;
// bram[5399] = 195;
// bram[5400] = 184;
// bram[5401] = 172;
// bram[5402] = 160;
// bram[5403] = 147;
// bram[5404] = 134;
// bram[5405] = 121;
// bram[5406] = 108;
// bram[5407] = 95;
// bram[5408] = 83;
// bram[5409] = 71;
// bram[5410] = 59;
// bram[5411] = 49;
// bram[5412] = 39;
// bram[5413] = 30;
// bram[5414] = 22;
// bram[5415] = 15;
// bram[5416] = 9;
// bram[5417] = 5;
// bram[5418] = 2;
// bram[5419] = 0;
// bram[5420] = 0;
// bram[5421] = 0;
// bram[5422] = 3;
// bram[5423] = 6;
// bram[5424] = 11;
// bram[5425] = 17;
// bram[5426] = 24;
// bram[5427] = 32;
// bram[5428] = 42;
// bram[5429] = 52;
// bram[5430] = 63;
// bram[5431] = 74;
// bram[5432] = 86;
// bram[5433] = 99;
// bram[5434] = 112;
// bram[5435] = 125;
// bram[5436] = 138;
// bram[5437] = 151;
// bram[5438] = 164;
// bram[5439] = 176;
// bram[5440] = 188;
// bram[5441] = 199;
// bram[5442] = 209;
// bram[5443] = 219;
// bram[5444] = 227;
// bram[5445] = 235;
// bram[5446] = 241;
// bram[5447] = 246;
// bram[5448] = 250;
// bram[5449] = 252;
// bram[5450] = 253;
// bram[5451] = 253;
// bram[5452] = 252;
// bram[5453] = 249;
// bram[5454] = 245;
// bram[5455] = 239;
// bram[5456] = 233;
// bram[5457] = 225;
// bram[5458] = 216;
// bram[5459] = 207;
// bram[5460] = 196;
// bram[5461] = 185;
// bram[5462] = 173;
// bram[5463] = 161;
// bram[5464] = 148;
// bram[5465] = 135;
// bram[5466] = 122;
// bram[5467] = 109;
// bram[5468] = 96;
// bram[5469] = 84;
// bram[5470] = 72;
// bram[5471] = 60;
// bram[5472] = 49;
// bram[5473] = 39;
// bram[5474] = 30;
// bram[5475] = 22;
// bram[5476] = 15;
// bram[5477] = 10;
// bram[5478] = 5;
// bram[5479] = 2;
// bram[5480] = 0;
// bram[5481] = 0;
// bram[5482] = 0;
// bram[5483] = 2;
// bram[5484] = 6;
// bram[5485] = 11;
// bram[5486] = 16;
// bram[5487] = 24;
// bram[5488] = 32;
// bram[5489] = 41;
// bram[5490] = 51;
// bram[5491] = 62;
// bram[5492] = 74;
// bram[5493] = 86;
// bram[5494] = 98;
// bram[5495] = 111;
// bram[5496] = 124;
// bram[5497] = 137;
// bram[5498] = 150;
// bram[5499] = 163;
// bram[5500] = 175;
// bram[5501] = 187;
// bram[5502] = 198;
// bram[5503] = 208;
// bram[5504] = 218;
// bram[5505] = 227;
// bram[5506] = 234;
// bram[5507] = 240;
// bram[5508] = 246;
// bram[5509] = 249;
// bram[5510] = 252;
// bram[5511] = 253;
// bram[5512] = 253;
// bram[5513] = 252;
// bram[5514] = 249;
// bram[5515] = 245;
// bram[5516] = 240;
// bram[5517] = 233;
// bram[5518] = 226;
// bram[5519] = 217;
// bram[5520] = 207;
// bram[5521] = 197;
// bram[5522] = 186;
// bram[5523] = 174;
// bram[5524] = 162;
// bram[5525] = 149;
// bram[5526] = 136;
// bram[5527] = 123;
// bram[5528] = 110;
// bram[5529] = 97;
// bram[5530] = 84;
// bram[5531] = 72;
// bram[5532] = 61;
// bram[5533] = 50;
// bram[5534] = 40;
// bram[5535] = 31;
// bram[5536] = 23;
// bram[5537] = 16;
// bram[5538] = 10;
// bram[5539] = 5;
// bram[5540] = 2;
// bram[5541] = 0;
// bram[5542] = 0;
// bram[5543] = 0;
// bram[5544] = 2;
// bram[5545] = 6;
// bram[5546] = 10;
// bram[5547] = 16;
// bram[5548] = 23;
// bram[5549] = 31;
// bram[5550] = 40;
// bram[5551] = 50;
// bram[5552] = 61;
// bram[5553] = 73;
// bram[5554] = 85;
// bram[5555] = 97;
// bram[5556] = 110;
// bram[5557] = 123;
// bram[5558] = 136;
// bram[5559] = 149;
// bram[5560] = 162;
// bram[5561] = 174;
// bram[5562] = 186;
// bram[5563] = 197;
// bram[5564] = 208;
// bram[5565] = 217;
// bram[5566] = 226;
// bram[5567] = 234;
// bram[5568] = 240;
// bram[5569] = 245;
// bram[5570] = 249;
// bram[5571] = 252;
// bram[5572] = 253;
// bram[5573] = 253;
// bram[5574] = 252;
// bram[5575] = 249;
// bram[5576] = 245;
// bram[5577] = 240;
// bram[5578] = 234;
// bram[5579] = 226;
// bram[5580] = 218;
// bram[5581] = 208;
// bram[5582] = 198;
// bram[5583] = 187;
// bram[5584] = 175;
// bram[5585] = 162;
// bram[5586] = 150;
// bram[5587] = 137;
// bram[5588] = 124;
// bram[5589] = 111;
// bram[5590] = 98;
// bram[5591] = 85;
// bram[5592] = 73;
// bram[5593] = 62;
// bram[5594] = 51;
// bram[5595] = 41;
// bram[5596] = 32;
// bram[5597] = 23;
// bram[5598] = 16;
// bram[5599] = 10;
// bram[5600] = 6;
// bram[5601] = 2;
// bram[5602] = 0;
// bram[5603] = 0;
// bram[5604] = 0;
// bram[5605] = 2;
// bram[5606] = 5;
// bram[5607] = 10;
// bram[5608] = 16;
// bram[5609] = 23;
// bram[5610] = 31;
// bram[5611] = 40;
// bram[5612] = 50;
// bram[5613] = 60;
// bram[5614] = 72;
// bram[5615] = 84;
// bram[5616] = 96;
// bram[5617] = 109;
// bram[5618] = 122;
// bram[5619] = 135;
// bram[5620] = 148;
// bram[5621] = 161;
// bram[5622] = 173;
// bram[5623] = 185;
// bram[5624] = 197;
// bram[5625] = 207;
// bram[5626] = 217;
// bram[5627] = 225;
// bram[5628] = 233;
// bram[5629] = 240;
// bram[5630] = 245;
// bram[5631] = 249;
// bram[5632] = 252;
// bram[5633] = 253;
// bram[5634] = 253;
// bram[5635] = 252;
// bram[5636] = 250;
// bram[5637] = 246;
// bram[5638] = 241;
// bram[5639] = 234;
// bram[5640] = 227;
// bram[5641] = 218;
// bram[5642] = 209;
// bram[5643] = 198;
// bram[5644] = 187;
// bram[5645] = 176;
// bram[5646] = 163;
// bram[5647] = 151;
// bram[5648] = 138;
// bram[5649] = 125;
// bram[5650] = 112;
// bram[5651] = 99;
// bram[5652] = 86;
// bram[5653] = 74;
// bram[5654] = 62;
// bram[5655] = 51;
// bram[5656] = 41;
// bram[5657] = 32;
// bram[5658] = 24;
// bram[5659] = 17;
// bram[5660] = 11;
// bram[5661] = 6;
// bram[5662] = 3;
// bram[5663] = 0;
// bram[5664] = 0;
// bram[5665] = 0;
// bram[5666] = 2;
// bram[5667] = 5;
// bram[5668] = 9;
// bram[5669] = 15;
// bram[5670] = 22;
// bram[5671] = 30;
// bram[5672] = 39;
// bram[5673] = 49;
// bram[5674] = 60;
// bram[5675] = 71;
// bram[5676] = 83;
// bram[5677] = 96;
// bram[5678] = 108;
// bram[5679] = 121;
// bram[5680] = 134;
// bram[5681] = 147;
// bram[5682] = 160;
// bram[5683] = 173;
// bram[5684] = 185;
// bram[5685] = 196;
// bram[5686] = 206;
// bram[5687] = 216;
// bram[5688] = 225;
// bram[5689] = 233;
// bram[5690] = 239;
// bram[5691] = 245;
// bram[5692] = 249;
// bram[5693] = 252;
// bram[5694] = 253;
// bram[5695] = 253;
// bram[5696] = 252;
// bram[5697] = 250;
// bram[5698] = 246;
// bram[5699] = 241;
// bram[5700] = 235;
// bram[5701] = 227;
// bram[5702] = 219;
// bram[5703] = 210;
// bram[5704] = 199;
// bram[5705] = 188;
// bram[5706] = 176;
// bram[5707] = 164;
// bram[5708] = 151;
// bram[5709] = 139;
// bram[5710] = 126;
// bram[5711] = 112;
// bram[5712] = 100;
// bram[5713] = 87;
// bram[5714] = 75;
// bram[5715] = 63;
// bram[5716] = 52;
// bram[5717] = 42;
// bram[5718] = 33;
// bram[5719] = 24;
// bram[5720] = 17;
// bram[5721] = 11;
// bram[5722] = 6;
// bram[5723] = 3;
// bram[5724] = 0;
// bram[5725] = 0;
// bram[5726] = 0;
// bram[5727] = 2;
// bram[5728] = 5;
// bram[5729] = 9;
// bram[5730] = 15;
// bram[5731] = 22;
// bram[5732] = 29;
// bram[5733] = 38;
// bram[5734] = 48;
// bram[5735] = 59;
// bram[5736] = 70;
// bram[5737] = 82;
// bram[5738] = 95;
// bram[5739] = 108;
// bram[5740] = 121;
// bram[5741] = 134;
// bram[5742] = 147;
// bram[5743] = 159;
// bram[5744] = 172;
// bram[5745] = 184;
// bram[5746] = 195;
// bram[5747] = 206;
// bram[5748] = 215;
// bram[5749] = 224;
// bram[5750] = 232;
// bram[5751] = 239;
// bram[5752] = 244;
// bram[5753] = 249;
// bram[5754] = 252;
// bram[5755] = 253;
// bram[5756] = 253;
// bram[5757] = 252;
// bram[5758] = 250;
// bram[5759] = 246;
// bram[5760] = 241;
// bram[5761] = 235;
// bram[5762] = 228;
// bram[5763] = 220;
// bram[5764] = 210;
// bram[5765] = 200;
// bram[5766] = 189;
// bram[5767] = 177;
// bram[5768] = 165;
// bram[5769] = 152;
// bram[5770] = 139;
// bram[5771] = 126;
// bram[5772] = 113;
// bram[5773] = 100;
// bram[5774] = 88;
// bram[5775] = 76;
// bram[5776] = 64;
// bram[5777] = 53;
// bram[5778] = 43;
// bram[5779] = 33;
// bram[5780] = 25;
// bram[5781] = 18;
// bram[5782] = 12;
// bram[5783] = 7;
// bram[5784] = 3;
// bram[5785] = 1;
// bram[5786] = 0;
// bram[5787] = 0;
// bram[5788] = 2;
// bram[5789] = 5;
// bram[5790] = 9;
// bram[5791] = 14;
// bram[5792] = 21;
// bram[5793] = 29;
// bram[5794] = 38;
// bram[5795] = 47;
// bram[5796] = 58;
// bram[5797] = 69;
// bram[5798] = 81;
// bram[5799] = 94;
// bram[5800] = 107;
// bram[5801] = 120;
// bram[5802] = 133;
// bram[5803] = 146;
// bram[5804] = 158;
// bram[5805] = 171;
// bram[5806] = 183;
// bram[5807] = 194;
// bram[5808] = 205;
// bram[5809] = 215;
// bram[5810] = 224;
// bram[5811] = 232;
// bram[5812] = 238;
// bram[5813] = 244;
// bram[5814] = 248;
// bram[5815] = 251;
// bram[5816] = 253;
// bram[5817] = 253;
// bram[5818] = 253;
// bram[5819] = 250;
// bram[5820] = 247;
// bram[5821] = 242;
// bram[5822] = 236;
// bram[5823] = 228;
// bram[5824] = 220;
// bram[5825] = 211;
// bram[5826] = 201;
// bram[5827] = 190;
// bram[5828] = 178;
// bram[5829] = 166;
// bram[5830] = 153;
// bram[5831] = 140;
// bram[5832] = 127;
// bram[5833] = 114;
// bram[5834] = 101;
// bram[5835] = 89;
// bram[5836] = 76;
// bram[5837] = 65;
// bram[5838] = 54;
// bram[5839] = 43;
// bram[5840] = 34;
// bram[5841] = 25;
// bram[5842] = 18;
// bram[5843] = 12;
// bram[5844] = 7;
// bram[5845] = 3;
// bram[5846] = 1;
// bram[5847] = 0;
// bram[5848] = 0;
// bram[5849] = 1;
// bram[5850] = 4;
// bram[5851] = 8;
// bram[5852] = 14;
// bram[5853] = 21;
// bram[5854] = 28;
// bram[5855] = 37;
// bram[5856] = 47;
// bram[5857] = 57;
// bram[5858] = 69;
// bram[5859] = 81;
// bram[5860] = 93;
// bram[5861] = 106;
// bram[5862] = 119;
// bram[5863] = 132;
// bram[5864] = 145;
// bram[5865] = 158;
// bram[5866] = 170;
// bram[5867] = 182;
// bram[5868] = 194;
// bram[5869] = 204;
// bram[5870] = 214;
// bram[5871] = 223;
// bram[5872] = 231;
// bram[5873] = 238;
// bram[5874] = 244;
// bram[5875] = 248;
// bram[5876] = 251;
// bram[5877] = 253;
// bram[5878] = 253;
// bram[5879] = 253;
// bram[5880] = 250;
// bram[5881] = 247;
// bram[5882] = 242;
// bram[5883] = 236;
// bram[5884] = 229;
// bram[5885] = 221;
// bram[5886] = 212;
// bram[5887] = 201;
// bram[5888] = 190;
// bram[5889] = 179;
// bram[5890] = 167;
// bram[5891] = 154;
// bram[5892] = 141;
// bram[5893] = 128;
// bram[5894] = 115;
// bram[5895] = 102;
// bram[5896] = 90;
// bram[5897] = 77;
// bram[5898] = 65;
// bram[5899] = 54;
// bram[5900] = 44;
// bram[5901] = 35;
// bram[5902] = 26;
// bram[5903] = 19;
// bram[5904] = 12;
// bram[5905] = 7;
// bram[5906] = 3;
// bram[5907] = 1;
// bram[5908] = 0;
// bram[5909] = 0;
// bram[5910] = 1;
// bram[5911] = 4;
// bram[5912] = 8;
// bram[5913] = 13;
// bram[5914] = 20;
// bram[5915] = 28;
// bram[5916] = 36;
// bram[5917] = 46;
// bram[5918] = 57;
// bram[5919] = 68;
// bram[5920] = 80;
// bram[5921] = 92;
// bram[5922] = 105;
// bram[5923] = 118;
// bram[5924] = 131;
// bram[5925] = 144;
// bram[5926] = 157;
// bram[5927] = 169;
// bram[5928] = 181;
// bram[5929] = 193;
// bram[5930] = 204;
// bram[5931] = 214;
// bram[5932] = 223;
// bram[5933] = 231;
// bram[5934] = 238;
// bram[5935] = 243;
// bram[5936] = 248;
// bram[5937] = 251;
// bram[5938] = 253;
// bram[5939] = 253;
// bram[5940] = 253;
// bram[5941] = 251;
// bram[5942] = 247;
// bram[5943] = 243;
// bram[5944] = 237;
// bram[5945] = 230;
// bram[5946] = 221;
// bram[5947] = 212;
// bram[5948] = 202;
// bram[5949] = 191;
// bram[5950] = 180;
// bram[5951] = 168;
// bram[5952] = 155;
// bram[5953] = 142;
// bram[5954] = 129;
// bram[5955] = 116;
// bram[5956] = 103;
// bram[5957] = 90;
// bram[5958] = 78;
// bram[5959] = 66;
// bram[5960] = 55;
// bram[5961] = 45;
// bram[5962] = 35;
// bram[5963] = 27;
// bram[5964] = 19;
// bram[5965] = 13;
// bram[5966] = 7;
// bram[5967] = 4;
// bram[5968] = 1;
// bram[5969] = 0;
// bram[5970] = 0;
// bram[5971] = 1;
// bram[5972] = 4;
// bram[5973] = 8;
// bram[5974] = 13;
// bram[5975] = 20;
// bram[5976] = 27;
// bram[5977] = 36;
// bram[5978] = 45;
// bram[5979] = 56;
// bram[5980] = 67;
// bram[5981] = 79;
// bram[5982] = 91;
// bram[5983] = 104;
// bram[5984] = 117;
// bram[5985] = 130;
// bram[5986] = 143;
// bram[5987] = 156;
// bram[5988] = 168;
// bram[5989] = 180;
// bram[5990] = 192;
// bram[5991] = 203;
// bram[5992] = 213;
// bram[5993] = 222;
// bram[5994] = 230;
// bram[5995] = 237;
// bram[5996] = 243;
// bram[5997] = 247;
// bram[5998] = 251;
// bram[5999] = 253;
// bram[6000] = 254;
// bram[6001] = 253;
// bram[6002] = 251;
// bram[6003] = 247;
// bram[6004] = 243;
// bram[6005] = 237;
// bram[6006] = 230;
// bram[6007] = 222;
// bram[6008] = 213;
// bram[6009] = 203;
// bram[6010] = 192;
// bram[6011] = 180;
// bram[6012] = 168;
// bram[6013] = 156;
// bram[6014] = 143;
// bram[6015] = 130;
// bram[6016] = 117;
// bram[6017] = 104;
// bram[6018] = 91;
// bram[6019] = 79;
// bram[6020] = 67;
// bram[6021] = 56;
// bram[6022] = 45;
// bram[6023] = 36;
// bram[6024] = 27;
// bram[6025] = 20;
// bram[6026] = 13;
// bram[6027] = 8;
// bram[6028] = 4;
// bram[6029] = 1;
// bram[6030] = 0;
// bram[6031] = 0;
// bram[6032] = 1;
// bram[6033] = 4;
// bram[6034] = 7;
// bram[6035] = 13;
// bram[6036] = 19;
// bram[6037] = 27;
// bram[6038] = 35;
// bram[6039] = 45;
// bram[6040] = 55;
// bram[6041] = 66;
// bram[6042] = 78;
// bram[6043] = 90;
// bram[6044] = 103;
// bram[6045] = 116;
// bram[6046] = 129;
// bram[6047] = 142;
// bram[6048] = 155;
// bram[6049] = 168;
// bram[6050] = 180;
// bram[6051] = 191;
// bram[6052] = 202;
// bram[6053] = 212;
// bram[6054] = 221;
// bram[6055] = 230;
// bram[6056] = 237;
// bram[6057] = 243;
// bram[6058] = 247;
// bram[6059] = 251;
// bram[6060] = 253;
// bram[6061] = 253;
// bram[6062] = 253;
// bram[6063] = 251;
// bram[6064] = 248;
// bram[6065] = 243;
// bram[6066] = 238;
// bram[6067] = 231;
// bram[6068] = 223;
// bram[6069] = 214;
// bram[6070] = 204;
// bram[6071] = 193;
// bram[6072] = 181;
// bram[6073] = 169;
// bram[6074] = 157;
// bram[6075] = 144;
// bram[6076] = 131;
// bram[6077] = 118;
// bram[6078] = 105;
// bram[6079] = 92;
// bram[6080] = 80;
// bram[6081] = 68;
// bram[6082] = 57;
// bram[6083] = 46;
// bram[6084] = 36;
// bram[6085] = 28;
// bram[6086] = 20;
// bram[6087] = 13;
// bram[6088] = 8;
// bram[6089] = 4;
// bram[6090] = 1;
// bram[6091] = 0;
// bram[6092] = 0;
// bram[6093] = 1;
// bram[6094] = 3;
// bram[6095] = 7;
// bram[6096] = 12;
// bram[6097] = 19;
// bram[6098] = 26;
// bram[6099] = 35;
// bram[6100] = 44;
// bram[6101] = 54;
// bram[6102] = 65;
// bram[6103] = 77;
// bram[6104] = 90;
// bram[6105] = 102;
// bram[6106] = 115;
// bram[6107] = 128;
// bram[6108] = 141;
// bram[6109] = 154;
// bram[6110] = 167;
// bram[6111] = 179;
// bram[6112] = 190;
// bram[6113] = 201;
// bram[6114] = 212;
// bram[6115] = 221;
// bram[6116] = 229;
// bram[6117] = 236;
// bram[6118] = 242;
// bram[6119] = 247;
// bram[6120] = 250;
// bram[6121] = 253;
// bram[6122] = 253;
// bram[6123] = 253;
// bram[6124] = 251;
// bram[6125] = 248;
// bram[6126] = 244;
// bram[6127] = 238;
// bram[6128] = 231;
// bram[6129] = 223;
// bram[6130] = 214;
// bram[6131] = 204;
// bram[6132] = 194;
// bram[6133] = 182;
// bram[6134] = 170;
// bram[6135] = 158;
// bram[6136] = 145;
// bram[6137] = 132;
// bram[6138] = 119;
// bram[6139] = 106;
// bram[6140] = 93;
// bram[6141] = 81;
// bram[6142] = 69;
// bram[6143] = 57;
// bram[6144] = 47;
// bram[6145] = 37;
// bram[6146] = 28;
// bram[6147] = 21;
// bram[6148] = 14;
// bram[6149] = 8;
// bram[6150] = 4;
// bram[6151] = 1;
// bram[6152] = 0;
// bram[6153] = 0;
// bram[6154] = 1;
// bram[6155] = 3;
// bram[6156] = 7;
// bram[6157] = 12;
// bram[6158] = 18;
// bram[6159] = 25;
// bram[6160] = 34;
// bram[6161] = 43;
// bram[6162] = 54;
// bram[6163] = 65;
// bram[6164] = 76;
// bram[6165] = 89;
// bram[6166] = 101;
// bram[6167] = 114;
// bram[6168] = 127;
// bram[6169] = 140;
// bram[6170] = 153;
// bram[6171] = 166;
// bram[6172] = 178;
// bram[6173] = 190;
// bram[6174] = 201;
// bram[6175] = 211;
// bram[6176] = 220;
// bram[6177] = 228;
// bram[6178] = 236;
// bram[6179] = 242;
// bram[6180] = 247;
// bram[6181] = 250;
// bram[6182] = 253;
// bram[6183] = 253;
// bram[6184] = 253;
// bram[6185] = 251;
// bram[6186] = 248;
// bram[6187] = 244;
// bram[6188] = 238;
// bram[6189] = 232;
// bram[6190] = 224;
// bram[6191] = 215;
// bram[6192] = 205;
// bram[6193] = 194;
// bram[6194] = 183;
// bram[6195] = 171;
// bram[6196] = 158;
// bram[6197] = 146;
// bram[6198] = 133;
// bram[6199] = 120;
// bram[6200] = 107;
// bram[6201] = 94;
// bram[6202] = 81;
// bram[6203] = 69;
// bram[6204] = 58;
// bram[6205] = 47;
// bram[6206] = 38;
// bram[6207] = 29;
// bram[6208] = 21;
// bram[6209] = 14;
// bram[6210] = 9;
// bram[6211] = 5;
// bram[6212] = 2;
// bram[6213] = 0;
// bram[6214] = 0;
// bram[6215] = 1;
// bram[6216] = 3;
// bram[6217] = 7;
// bram[6218] = 12;
// bram[6219] = 18;
// bram[6220] = 25;
// bram[6221] = 33;
// bram[6222] = 43;
// bram[6223] = 53;
// bram[6224] = 64;
// bram[6225] = 76;
// bram[6226] = 88;
// bram[6227] = 100;
// bram[6228] = 113;
// bram[6229] = 126;
// bram[6230] = 139;
// bram[6231] = 152;
// bram[6232] = 165;
// bram[6233] = 177;
// bram[6234] = 189;
// bram[6235] = 200;
// bram[6236] = 210;
// bram[6237] = 220;
// bram[6238] = 228;
// bram[6239] = 235;
// bram[6240] = 241;
// bram[6241] = 246;
// bram[6242] = 250;
// bram[6243] = 252;
// bram[6244] = 253;
// bram[6245] = 253;
// bram[6246] = 252;
// bram[6247] = 249;
// bram[6248] = 244;
// bram[6249] = 239;
// bram[6250] = 232;
// bram[6251] = 224;
// bram[6252] = 215;
// bram[6253] = 206;
// bram[6254] = 195;
// bram[6255] = 184;
// bram[6256] = 172;
// bram[6257] = 159;
// bram[6258] = 147;
// bram[6259] = 134;
// bram[6260] = 121;
// bram[6261] = 108;
// bram[6262] = 95;
// bram[6263] = 82;
// bram[6264] = 70;
// bram[6265] = 59;
// bram[6266] = 48;
// bram[6267] = 38;
// bram[6268] = 29;
// bram[6269] = 22;
// bram[6270] = 15;
// bram[6271] = 9;
// bram[6272] = 5;
// bram[6273] = 2;
// bram[6274] = 0;
// bram[6275] = 0;
// bram[6276] = 0;
// bram[6277] = 3;
// bram[6278] = 6;
// bram[6279] = 11;
// bram[6280] = 17;
// bram[6281] = 24;
// bram[6282] = 33;
// bram[6283] = 42;
// bram[6284] = 52;
// bram[6285] = 63;
// bram[6286] = 75;
// bram[6287] = 87;
// bram[6288] = 100;
// bram[6289] = 112;
// bram[6290] = 126;
// bram[6291] = 139;
// bram[6292] = 151;
// bram[6293] = 164;
// bram[6294] = 176;
// bram[6295] = 188;
// bram[6296] = 199;
// bram[6297] = 210;
// bram[6298] = 219;
// bram[6299] = 227;
// bram[6300] = 235;
// bram[6301] = 241;
// bram[6302] = 246;
// bram[6303] = 250;
// bram[6304] = 252;
// bram[6305] = 253;
// bram[6306] = 253;
// bram[6307] = 252;
// bram[6308] = 249;
// bram[6309] = 245;
// bram[6310] = 239;
// bram[6311] = 233;
// bram[6312] = 225;
// bram[6313] = 216;
// bram[6314] = 206;
// bram[6315] = 196;
// bram[6316] = 185;
// bram[6317] = 173;
// bram[6318] = 160;
// bram[6319] = 147;
// bram[6320] = 134;
// bram[6321] = 121;
// bram[6322] = 108;
// bram[6323] = 96;
// bram[6324] = 83;
// bram[6325] = 71;
// bram[6326] = 60;
// bram[6327] = 49;
// bram[6328] = 39;
// bram[6329] = 30;
// bram[6330] = 22;
// bram[6331] = 15;
// bram[6332] = 9;
// bram[6333] = 5;
// bram[6334] = 2;
// bram[6335] = 0;
// bram[6336] = 0;
// bram[6337] = 0;
// bram[6338] = 3;
// bram[6339] = 6;
// bram[6340] = 11;
// bram[6341] = 17;
// bram[6342] = 24;
// bram[6343] = 32;
// bram[6344] = 41;
// bram[6345] = 51;
// bram[6346] = 62;
// bram[6347] = 74;
// bram[6348] = 86;
// bram[6349] = 99;
// bram[6350] = 112;
// bram[6351] = 125;
// bram[6352] = 138;
// bram[6353] = 151;
// bram[6354] = 163;
// bram[6355] = 176;
// bram[6356] = 187;
// bram[6357] = 198;
// bram[6358] = 209;
// bram[6359] = 218;
// bram[6360] = 227;
// bram[6361] = 234;
// bram[6362] = 241;
// bram[6363] = 246;
// bram[6364] = 250;
// bram[6365] = 252;
// bram[6366] = 253;
// bram[6367] = 253;
// bram[6368] = 252;
// bram[6369] = 249;
// bram[6370] = 245;
// bram[6371] = 240;
// bram[6372] = 233;
// bram[6373] = 225;
// bram[6374] = 217;
// bram[6375] = 207;
// bram[6376] = 197;
// bram[6377] = 185;
// bram[6378] = 173;
// bram[6379] = 161;
// bram[6380] = 148;
// bram[6381] = 135;
// bram[6382] = 122;
// bram[6383] = 109;
// bram[6384] = 96;
// bram[6385] = 84;
// bram[6386] = 72;
// bram[6387] = 60;
// bram[6388] = 50;
// bram[6389] = 40;
// bram[6390] = 31;
// bram[6391] = 23;
// bram[6392] = 16;
// bram[6393] = 10;
// bram[6394] = 5;
// bram[6395] = 2;
// bram[6396] = 0;
// bram[6397] = 0;
// bram[6398] = 0;
// bram[6399] = 2;
// bram[6400] = 6;
// bram[6401] = 10;
// bram[6402] = 16;
// bram[6403] = 23;
// bram[6404] = 32;
// bram[6405] = 41;
// bram[6406] = 51;
// bram[6407] = 62;
// bram[6408] = 73;
// bram[6409] = 85;
// bram[6410] = 98;
// bram[6411] = 111;
// bram[6412] = 124;
// bram[6413] = 137;
// bram[6414] = 150;
// bram[6415] = 162;
// bram[6416] = 175;
// bram[6417] = 187;
// bram[6418] = 198;
// bram[6419] = 208;
// bram[6420] = 218;
// bram[6421] = 226;
// bram[6422] = 234;
// bram[6423] = 240;
// bram[6424] = 245;
// bram[6425] = 249;
// bram[6426] = 252;
// bram[6427] = 253;
// bram[6428] = 253;
// bram[6429] = 252;
// bram[6430] = 249;
// bram[6431] = 245;
// bram[6432] = 240;
// bram[6433] = 234;
// bram[6434] = 226;
// bram[6435] = 217;
// bram[6436] = 208;
// bram[6437] = 197;
// bram[6438] = 186;
// bram[6439] = 174;
// bram[6440] = 162;
// bram[6441] = 149;
// bram[6442] = 136;
// bram[6443] = 123;
// bram[6444] = 110;
// bram[6445] = 97;
// bram[6446] = 85;
// bram[6447] = 73;
// bram[6448] = 61;
// bram[6449] = 50;
// bram[6450] = 40;
// bram[6451] = 31;
// bram[6452] = 23;
// bram[6453] = 16;
// bram[6454] = 10;
// bram[6455] = 6;
// bram[6456] = 2;
// bram[6457] = 0;
// bram[6458] = 0;
// bram[6459] = 0;
// bram[6460] = 2;
// bram[6461] = 5;
// bram[6462] = 10;
// bram[6463] = 16;
// bram[6464] = 23;
// bram[6465] = 31;
// bram[6466] = 40;
// bram[6467] = 50;
// bram[6468] = 61;
// bram[6469] = 72;
// bram[6470] = 84;
// bram[6471] = 97;
// bram[6472] = 110;
// bram[6473] = 123;
// bram[6474] = 136;
// bram[6475] = 149;
// bram[6476] = 162;
// bram[6477] = 174;
// bram[6478] = 186;
// bram[6479] = 197;
// bram[6480] = 207;
// bram[6481] = 217;
// bram[6482] = 226;
// bram[6483] = 233;
// bram[6484] = 240;
// bram[6485] = 245;
// bram[6486] = 249;
// bram[6487] = 252;
// bram[6488] = 253;
// bram[6489] = 253;
// bram[6490] = 252;
// bram[6491] = 249;
// bram[6492] = 246;
// bram[6493] = 240;
// bram[6494] = 234;
// bram[6495] = 227;
// bram[6496] = 218;
// bram[6497] = 208;
// bram[6498] = 198;
// bram[6499] = 187;
// bram[6500] = 175;
// bram[6501] = 163;
// bram[6502] = 150;
// bram[6503] = 137;
// bram[6504] = 124;
// bram[6505] = 111;
// bram[6506] = 98;
// bram[6507] = 86;
// bram[6508] = 74;
// bram[6509] = 62;
// bram[6510] = 51;
// bram[6511] = 41;
// bram[6512] = 32;
// bram[6513] = 24;
// bram[6514] = 16;
// bram[6515] = 11;
// bram[6516] = 6;
// bram[6517] = 2;
// bram[6518] = 0;
// bram[6519] = 0;
// bram[6520] = 0;
// bram[6521] = 2;
// bram[6522] = 5;
// bram[6523] = 10;
// bram[6524] = 15;
// bram[6525] = 22;
// bram[6526] = 30;
// bram[6527] = 39;
// bram[6528] = 49;
// bram[6529] = 60;
// bram[6530] = 72;
// bram[6531] = 84;
// bram[6532] = 96;
// bram[6533] = 109;
// bram[6534] = 122;
// bram[6535] = 135;
// bram[6536] = 148;
// bram[6537] = 161;
// bram[6538] = 173;
// bram[6539] = 185;
// bram[6540] = 196;
// bram[6541] = 207;
// bram[6542] = 216;
// bram[6543] = 225;
// bram[6544] = 233;
// bram[6545] = 239;
// bram[6546] = 245;
// bram[6547] = 249;
// bram[6548] = 252;
// bram[6549] = 253;
// bram[6550] = 253;
// bram[6551] = 252;
// bram[6552] = 250;
// bram[6553] = 246;
// bram[6554] = 241;
// bram[6555] = 235;
// bram[6556] = 227;
// bram[6557] = 219;
// bram[6558] = 209;
// bram[6559] = 199;
// bram[6560] = 188;
// bram[6561] = 176;
// bram[6562] = 164;
// bram[6563] = 151;
// bram[6564] = 138;
// bram[6565] = 125;
// bram[6566] = 112;
// bram[6567] = 99;
// bram[6568] = 86;
// bram[6569] = 74;
// bram[6570] = 63;
// bram[6571] = 52;
// bram[6572] = 42;
// bram[6573] = 32;
// bram[6574] = 24;
// bram[6575] = 17;
// bram[6576] = 11;
// bram[6577] = 6;
// bram[6578] = 3;
// bram[6579] = 0;
// bram[6580] = 0;
// bram[6581] = 0;
// bram[6582] = 2;
// bram[6583] = 5;
// bram[6584] = 9;
// bram[6585] = 15;
// bram[6586] = 22;
// bram[6587] = 30;
// bram[6588] = 39;
// bram[6589] = 49;
// bram[6590] = 59;
// bram[6591] = 71;
// bram[6592] = 83;
// bram[6593] = 95;
// bram[6594] = 108;
// bram[6595] = 121;
// bram[6596] = 134;
// bram[6597] = 147;
// bram[6598] = 160;
// bram[6599] = 172;
// bram[6600] = 184;
// bram[6601] = 195;
// bram[6602] = 206;
// bram[6603] = 216;
// bram[6604] = 225;
// bram[6605] = 232;
// bram[6606] = 239;
// bram[6607] = 244;
// bram[6608] = 249;
// bram[6609] = 252;
// bram[6610] = 253;
// bram[6611] = 253;
// bram[6612] = 252;
// bram[6613] = 250;
// bram[6614] = 246;
// bram[6615] = 241;
// bram[6616] = 235;
// bram[6617] = 228;
// bram[6618] = 219;
// bram[6619] = 210;
// bram[6620] = 200;
// bram[6621] = 188;
// bram[6622] = 177;
// bram[6623] = 165;
// bram[6624] = 152;
// bram[6625] = 139;
// bram[6626] = 126;
// bram[6627] = 113;
// bram[6628] = 100;
// bram[6629] = 87;
// bram[6630] = 75;
// bram[6631] = 63;
// bram[6632] = 52;
// bram[6633] = 42;
// bram[6634] = 33;
// bram[6635] = 25;
// bram[6636] = 17;
// bram[6637] = 11;
// bram[6638] = 6;
// bram[6639] = 3;
// bram[6640] = 1;
// bram[6641] = 0;
// bram[6642] = 0;
// bram[6643] = 2;
// bram[6644] = 5;
// bram[6645] = 9;
// bram[6646] = 15;
// bram[6647] = 21;
// bram[6648] = 29;
// bram[6649] = 38;
// bram[6650] = 48;
// bram[6651] = 59;
// bram[6652] = 70;
// bram[6653] = 82;
// bram[6654] = 94;
// bram[6655] = 107;
// bram[6656] = 120;
// bram[6657] = 133;
// bram[6658] = 146;
// bram[6659] = 159;
// bram[6660] = 171;
// bram[6661] = 183;
// bram[6662] = 195;
// bram[6663] = 205;
// bram[6664] = 215;
// bram[6665] = 224;
// bram[6666] = 232;
// bram[6667] = 239;
// bram[6668] = 244;
// bram[6669] = 248;
// bram[6670] = 251;
// bram[6671] = 253;
// bram[6672] = 253;
// bram[6673] = 252;
// bram[6674] = 250;
// bram[6675] = 246;
// bram[6676] = 242;
// bram[6677] = 235;
// bram[6678] = 228;
// bram[6679] = 220;
// bram[6680] = 210;
// bram[6681] = 200;
// bram[6682] = 189;
// bram[6683] = 178;
// bram[6684] = 165;
// bram[6685] = 153;
// bram[6686] = 140;
// bram[6687] = 127;
// bram[6688] = 114;
// bram[6689] = 101;
// bram[6690] = 88;
// bram[6691] = 76;
// bram[6692] = 64;
// bram[6693] = 53;
// bram[6694] = 43;
// bram[6695] = 34;
// bram[6696] = 25;
// bram[6697] = 18;
// bram[6698] = 12;
// bram[6699] = 7;
// bram[6700] = 3;
// bram[6701] = 1;
// bram[6702] = 0;
// bram[6703] = 0;
// bram[6704] = 1;
// bram[6705] = 4;
// bram[6706] = 9;
// bram[6707] = 14;
// bram[6708] = 21;
// bram[6709] = 29;
// bram[6710] = 37;
// bram[6711] = 47;
// bram[6712] = 58;
// bram[6713] = 69;
// bram[6714] = 81;
// bram[6715] = 93;
// bram[6716] = 106;
// bram[6717] = 119;
// bram[6718] = 132;
// bram[6719] = 145;
// bram[6720] = 158;
// bram[6721] = 171;
// bram[6722] = 183;
// bram[6723] = 194;
// bram[6724] = 205;
// bram[6725] = 215;
// bram[6726] = 223;
// bram[6727] = 231;
// bram[6728] = 238;
// bram[6729] = 244;
// bram[6730] = 248;
// bram[6731] = 251;
// bram[6732] = 253;
// bram[6733] = 253;
// bram[6734] = 253;
// bram[6735] = 250;
// bram[6736] = 247;
// bram[6737] = 242;
// bram[6738] = 236;
// bram[6739] = 229;
// bram[6740] = 220;
// bram[6741] = 211;
// bram[6742] = 201;
// bram[6743] = 190;
// bram[6744] = 178;
// bram[6745] = 166;
// bram[6746] = 154;
// bram[6747] = 141;
// bram[6748] = 128;
// bram[6749] = 115;
// bram[6750] = 102;
// bram[6751] = 89;
// bram[6752] = 77;
// bram[6753] = 65;
// bram[6754] = 54;
// bram[6755] = 44;
// bram[6756] = 34;
// bram[6757] = 26;
// bram[6758] = 18;
// bram[6759] = 12;
// bram[6760] = 7;
// bram[6761] = 3;
// bram[6762] = 1;
// bram[6763] = 0;
// bram[6764] = 0;
// bram[6765] = 1;
// bram[6766] = 4;
// bram[6767] = 8;
// bram[6768] = 14;
// bram[6769] = 20;
// bram[6770] = 28;
// bram[6771] = 37;
// bram[6772] = 46;
// bram[6773] = 57;
// bram[6774] = 68;
// bram[6775] = 80;
// bram[6776] = 93;
// bram[6777] = 105;
// bram[6778] = 118;
// bram[6779] = 131;
// bram[6780] = 144;
// bram[6781] = 157;
// bram[6782] = 170;
// bram[6783] = 182;
// bram[6784] = 193;
// bram[6785] = 204;
// bram[6786] = 214;
// bram[6787] = 223;
// bram[6788] = 231;
// bram[6789] = 238;
// bram[6790] = 243;
// bram[6791] = 248;
// bram[6792] = 251;
// bram[6793] = 253;
// bram[6794] = 253;
// bram[6795] = 253;
// bram[6796] = 251;
// bram[6797] = 247;
// bram[6798] = 242;
// bram[6799] = 236;
// bram[6800] = 229;
// bram[6801] = 221;
// bram[6802] = 212;
// bram[6803] = 202;
// bram[6804] = 191;
// bram[6805] = 179;
// bram[6806] = 167;
// bram[6807] = 154;
// bram[6808] = 142;
// bram[6809] = 129;
// bram[6810] = 116;
// bram[6811] = 103;
// bram[6812] = 90;
// bram[6813] = 78;
// bram[6814] = 66;
// bram[6815] = 55;
// bram[6816] = 44;
// bram[6817] = 35;
// bram[6818] = 26;
// bram[6819] = 19;
// bram[6820] = 12;
// bram[6821] = 7;
// bram[6822] = 3;
// bram[6823] = 1;
// bram[6824] = 0;
// bram[6825] = 0;
// bram[6826] = 1;
// bram[6827] = 4;
// bram[6828] = 8;
// bram[6829] = 13;
// bram[6830] = 20;
// bram[6831] = 27;
// bram[6832] = 36;
// bram[6833] = 46;
// bram[6834] = 56;
// bram[6835] = 68;
// bram[6836] = 79;
// bram[6837] = 92;
// bram[6838] = 104;
// bram[6839] = 117;
// bram[6840] = 130;
// bram[6841] = 144;
// bram[6842] = 156;
// bram[6843] = 169;
// bram[6844] = 181;
// bram[6845] = 192;
// bram[6846] = 203;
// bram[6847] = 213;
// bram[6848] = 222;
// bram[6849] = 230;
// bram[6850] = 237;
// bram[6851] = 243;
// bram[6852] = 248;
// bram[6853] = 251;
// bram[6854] = 253;
// bram[6855] = 253;
// bram[6856] = 253;
// bram[6857] = 251;
// bram[6858] = 247;
// bram[6859] = 243;
// bram[6860] = 237;
// bram[6861] = 230;
// bram[6862] = 222;
// bram[6863] = 212;
// bram[6864] = 202;
// bram[6865] = 192;
// bram[6866] = 180;
// bram[6867] = 168;
// bram[6868] = 155;
// bram[6869] = 143;
// bram[6870] = 129;
// bram[6871] = 116;
// bram[6872] = 103;
// bram[6873] = 91;
// bram[6874] = 78;
// bram[6875] = 67;
// bram[6876] = 55;
// bram[6877] = 45;
// bram[6878] = 35;
// bram[6879] = 27;
// bram[6880] = 19;
// bram[6881] = 13;
// bram[6882] = 8;
// bram[6883] = 4;
// bram[6884] = 1;
// bram[6885] = 0;
// bram[6886] = 0;
// bram[6887] = 1;
// bram[6888] = 4;
// bram[6889] = 8;
// bram[6890] = 13;
// bram[6891] = 19;
// bram[6892] = 27;
// bram[6893] = 36;
// bram[6894] = 45;
// bram[6895] = 56;
// bram[6896] = 67;
// bram[6897] = 79;
// bram[6898] = 91;
// bram[6899] = 104;
// bram[6900] = 117;
// bram[6901] = 130;
// bram[6902] = 143;
// bram[6903] = 155;
// bram[6904] = 168;
// bram[6905] = 180;
// bram[6906] = 192;
// bram[6907] = 203;
// bram[6908] = 213;
// bram[6909] = 222;
// bram[6910] = 230;
// bram[6911] = 237;
// bram[6912] = 243;
// bram[6913] = 247;
// bram[6914] = 251;
// bram[6915] = 253;
// bram[6916] = 253;
// bram[6917] = 253;
// bram[6918] = 251;
// bram[6919] = 248;
// bram[6920] = 243;
// bram[6921] = 237;
// bram[6922] = 230;
// bram[6923] = 222;
// bram[6924] = 213;
// bram[6925] = 203;
// bram[6926] = 192;
// bram[6927] = 181;
// bram[6928] = 169;
// bram[6929] = 156;
// bram[6930] = 143;
// bram[6931] = 130;
// bram[6932] = 117;
// bram[6933] = 104;
// bram[6934] = 92;
// bram[6935] = 79;
// bram[6936] = 67;
// bram[6937] = 56;
// bram[6938] = 46;
// bram[6939] = 36;
// bram[6940] = 27;
// bram[6941] = 20;
// bram[6942] = 13;
// bram[6943] = 8;
// bram[6944] = 4;
// bram[6945] = 1;
// bram[6946] = 0;
// bram[6947] = 0;
// bram[6948] = 1;
// bram[6949] = 3;
// bram[6950] = 7;
// bram[6951] = 12;
// bram[6952] = 19;
// bram[6953] = 26;
// bram[6954] = 35;
// bram[6955] = 44;
// bram[6956] = 55;
// bram[6957] = 66;
// bram[6958] = 78;
// bram[6959] = 90;
// bram[6960] = 103;
// bram[6961] = 116;
// bram[6962] = 129;
// bram[6963] = 142;
// bram[6964] = 155;
// bram[6965] = 167;
// bram[6966] = 179;
// bram[6967] = 191;
// bram[6968] = 202;
// bram[6969] = 212;
// bram[6970] = 221;
// bram[6971] = 229;
// bram[6972] = 236;
// bram[6973] = 242;
// bram[6974] = 247;
// bram[6975] = 251;
// bram[6976] = 253;
// bram[6977] = 253;
// bram[6978] = 253;
// bram[6979] = 251;
// bram[6980] = 248;
// bram[6981] = 243;
// bram[6982] = 238;
// bram[6983] = 231;
// bram[6984] = 223;
// bram[6985] = 214;
// bram[6986] = 204;
// bram[6987] = 193;
// bram[6988] = 182;
// bram[6989] = 170;
// bram[6990] = 157;
// bram[6991] = 144;
// bram[6992] = 131;
// bram[6993] = 118;
// bram[6994] = 105;
// bram[6995] = 93;
// bram[6996] = 80;
// bram[6997] = 68;
// bram[6998] = 57;
// bram[6999] = 46;
// bram[7000] = 37;
// bram[7001] = 28;
// bram[7002] = 20;
// bram[7003] = 14;
// bram[7004] = 8;
// bram[7005] = 4;
// bram[7006] = 1;
// bram[7007] = 0;
// bram[7008] = 0;
// bram[7009] = 1;
// bram[7010] = 3;
// bram[7011] = 7;
// bram[7012] = 12;
// bram[7013] = 18;
// bram[7014] = 26;
// bram[7015] = 34;
// bram[7016] = 44;
// bram[7017] = 54;
// bram[7018] = 65;
// bram[7019] = 77;
// bram[7020] = 89;
// bram[7021] = 102;
// bram[7022] = 115;
// bram[7023] = 128;
// bram[7024] = 141;
// bram[7025] = 154;
// bram[7026] = 166;
// bram[7027] = 178;
// bram[7028] = 190;
// bram[7029] = 201;
// bram[7030] = 211;
// bram[7031] = 221;
// bram[7032] = 229;
// bram[7033] = 236;
// bram[7034] = 242;
// bram[7035] = 247;
// bram[7036] = 250;
// bram[7037] = 253;
// bram[7038] = 253;
// bram[7039] = 253;
// bram[7040] = 251;
// bram[7041] = 248;
// bram[7042] = 244;
// bram[7043] = 238;
// bram[7044] = 231;
// bram[7045] = 223;
// bram[7046] = 214;
// bram[7047] = 205;
// bram[7048] = 194;
// bram[7049] = 182;
// bram[7050] = 170;
// bram[7051] = 158;
// bram[7052] = 145;
// bram[7053] = 132;
// bram[7054] = 119;
// bram[7055] = 106;
// bram[7056] = 93;
// bram[7057] = 81;
// bram[7058] = 69;
// bram[7059] = 58;
// bram[7060] = 47;
// bram[7061] = 37;
// bram[7062] = 29;
// bram[7063] = 21;
// bram[7064] = 14;
// bram[7065] = 9;
// bram[7066] = 4;
// bram[7067] = 1;
// bram[7068] = 0;
// bram[7069] = 0;
// bram[7070] = 1;
// bram[7071] = 3;
// bram[7072] = 7;
// bram[7073] = 12;
// bram[7074] = 18;
// bram[7075] = 25;
// bram[7076] = 34;
// bram[7077] = 43;
// bram[7078] = 53;
// bram[7079] = 64;
// bram[7080] = 76;
// bram[7081] = 88;
// bram[7082] = 101;
// bram[7083] = 114;
// bram[7084] = 127;
// bram[7085] = 140;
// bram[7086] = 153;
// bram[7087] = 165;
// bram[7088] = 178;
// bram[7089] = 189;
// bram[7090] = 200;
// bram[7091] = 211;
// bram[7092] = 220;
// bram[7093] = 228;
// bram[7094] = 236;
// bram[7095] = 242;
// bram[7096] = 247;
// bram[7097] = 250;
// bram[7098] = 252;
// bram[7099] = 253;
// bram[7100] = 253;
// bram[7101] = 251;
// bram[7102] = 248;
// bram[7103] = 244;
// bram[7104] = 239;
// bram[7105] = 232;
// bram[7106] = 224;
// bram[7107] = 215;
// bram[7108] = 205;
// bram[7109] = 195;
// bram[7110] = 183;
// bram[7111] = 171;
// bram[7112] = 159;
// bram[7113] = 146;
// bram[7114] = 133;
// bram[7115] = 120;
// bram[7116] = 107;
// bram[7117] = 94;
// bram[7118] = 82;
// bram[7119] = 70;
// bram[7120] = 58;
// bram[7121] = 48;
// bram[7122] = 38;
// bram[7123] = 29;
// bram[7124] = 21;
// bram[7125] = 14;
// bram[7126] = 9;
// bram[7127] = 5;
// bram[7128] = 2;
// bram[7129] = 0;
// bram[7130] = 0;
// bram[7131] = 1;
// bram[7132] = 3;
// bram[7133] = 6;
// bram[7134] = 11;
// bram[7135] = 17;
// bram[7136] = 25;
// bram[7137] = 33;
// bram[7138] = 42;
// bram[7139] = 53;
// bram[7140] = 64;
// bram[7141] = 75;
// bram[7142] = 87;
// bram[7143] = 100;
// bram[7144] = 113;
// bram[7145] = 126;
// bram[7146] = 139;
// bram[7147] = 152;
// bram[7148] = 165;
// bram[7149] = 177;
// bram[7150] = 189;
// bram[7151] = 200;
// bram[7152] = 210;
// bram[7153] = 219;
// bram[7154] = 228;
// bram[7155] = 235;
// bram[7156] = 241;
// bram[7157] = 246;
// bram[7158] = 250;
// bram[7159] = 252;
// bram[7160] = 253;
// bram[7161] = 253;
// bram[7162] = 252;
// bram[7163] = 249;
// bram[7164] = 244;
// bram[7165] = 239;
// bram[7166] = 232;
// bram[7167] = 225;
// bram[7168] = 216;
// bram[7169] = 206;
// bram[7170] = 195;
// bram[7171] = 184;
// bram[7172] = 172;
// bram[7173] = 160;
// bram[7174] = 147;
// bram[7175] = 134;
// bram[7176] = 121;
// bram[7177] = 108;
// bram[7178] = 95;
// bram[7179] = 83;
// bram[7180] = 71;
// bram[7181] = 59;
// bram[7182] = 49;
// bram[7183] = 39;
// bram[7184] = 30;
// bram[7185] = 22;
// bram[7186] = 15;
// bram[7187] = 9;
// bram[7188] = 5;
// bram[7189] = 2;
// bram[7190] = 0;
// bram[7191] = 0;
// bram[7192] = 0;
// bram[7193] = 3;
// bram[7194] = 6;
// bram[7195] = 11;
// bram[7196] = 17;
// bram[7197] = 24;
// bram[7198] = 32;
// bram[7199] = 42;
// bram[7200] = 52;
// bram[7201] = 63;
// bram[7202] = 74;
// bram[7203] = 87;
// bram[7204] = 99;
// bram[7205] = 112;
// bram[7206] = 125;
// bram[7207] = 138;
// bram[7208] = 151;
// bram[7209] = 164;
// bram[7210] = 176;
// bram[7211] = 188;
// bram[7212] = 199;
// bram[7213] = 209;
// bram[7214] = 219;
// bram[7215] = 227;
// bram[7216] = 235;
// bram[7217] = 241;
// bram[7218] = 246;
// bram[7219] = 250;
// bram[7220] = 252;
// bram[7221] = 253;
// bram[7222] = 253;
// bram[7223] = 252;
// bram[7224] = 249;
// bram[7225] = 245;
// bram[7226] = 239;
// bram[7227] = 233;
// bram[7228] = 225;
// bram[7229] = 216;
// bram[7230] = 207;
// bram[7231] = 196;
// bram[7232] = 185;
// bram[7233] = 173;
// bram[7234] = 161;
// bram[7235] = 148;
// bram[7236] = 135;
// bram[7237] = 122;
// bram[7238] = 109;
// bram[7239] = 96;
// bram[7240] = 83;
// bram[7241] = 71;
// bram[7242] = 60;
// bram[7243] = 49;
// bram[7244] = 39;
// bram[7245] = 30;
// bram[7246] = 22;
// bram[7247] = 15;
// bram[7248] = 10;
// bram[7249] = 5;
// bram[7250] = 2;
// bram[7251] = 0;
// bram[7252] = 0;
// bram[7253] = 0;
// bram[7254] = 2;
// bram[7255] = 6;
// bram[7256] = 11;
// bram[7257] = 17;
// bram[7258] = 24;
// bram[7259] = 32;
// bram[7260] = 41;
// bram[7261] = 51;
// bram[7262] = 62;
// bram[7263] = 74;
// bram[7264] = 86;
// bram[7265] = 98;
// bram[7266] = 111;
// bram[7267] = 124;
// bram[7268] = 137;
// bram[7269] = 150;
// bram[7270] = 163;
// bram[7271] = 175;
// bram[7272] = 187;
// bram[7273] = 198;
// bram[7274] = 209;
// bram[7275] = 218;
// bram[7276] = 227;
// bram[7277] = 234;
// bram[7278] = 240;
// bram[7279] = 246;
// bram[7280] = 250;
// bram[7281] = 252;
// bram[7282] = 253;
// bram[7283] = 253;
// bram[7284] = 252;
// bram[7285] = 249;
// bram[7286] = 245;
// bram[7287] = 240;
// bram[7288] = 233;
// bram[7289] = 226;
// bram[7290] = 217;
// bram[7291] = 207;
// bram[7292] = 197;
// bram[7293] = 186;
// bram[7294] = 174;
// bram[7295] = 161;
// bram[7296] = 149;
// bram[7297] = 136;
// bram[7298] = 123;
// bram[7299] = 110;
// bram[7300] = 97;
// bram[7301] = 84;
// bram[7302] = 72;
// bram[7303] = 61;
// bram[7304] = 50;
// bram[7305] = 40;
// bram[7306] = 31;
// bram[7307] = 23;
// bram[7308] = 16;
// bram[7309] = 10;
// bram[7310] = 5;
// bram[7311] = 2;
// bram[7312] = 0;
// bram[7313] = 0;
// bram[7314] = 0;
// bram[7315] = 2;
// bram[7316] = 6;
// bram[7317] = 10;
// bram[7318] = 16;
// bram[7319] = 23;
// bram[7320] = 31;
// bram[7321] = 40;
// bram[7322] = 50;
// bram[7323] = 61;
// bram[7324] = 73;
// bram[7325] = 85;
// bram[7326] = 97;
// bram[7327] = 110;
// bram[7328] = 123;
// bram[7329] = 136;
// bram[7330] = 149;
// bram[7331] = 162;
// bram[7332] = 174;
// bram[7333] = 186;
// bram[7334] = 197;
// bram[7335] = 208;
// bram[7336] = 217;
// bram[7337] = 226;
// bram[7338] = 234;
// bram[7339] = 240;
// bram[7340] = 245;
// bram[7341] = 249;
// bram[7342] = 252;
// bram[7343] = 253;
// bram[7344] = 253;
// bram[7345] = 252;
// bram[7346] = 249;
// bram[7347] = 245;
// bram[7348] = 240;
// bram[7349] = 234;
// bram[7350] = 226;
// bram[7351] = 218;
// bram[7352] = 208;
// bram[7353] = 198;
// bram[7354] = 186;
// bram[7355] = 175;
// bram[7356] = 162;
// bram[7357] = 150;
// bram[7358] = 137;
// bram[7359] = 124;
// bram[7360] = 111;
// bram[7361] = 98;
// bram[7362] = 85;
// bram[7363] = 73;
// bram[7364] = 62;
// bram[7365] = 51;
// bram[7366] = 41;
// bram[7367] = 31;
// bram[7368] = 23;
// bram[7369] = 16;
// bram[7370] = 10;
// bram[7371] = 6;
// bram[7372] = 2;
// bram[7373] = 0;
// bram[7374] = 0;
// bram[7375] = 0;
// bram[7376] = 2;
// bram[7377] = 5;
// bram[7378] = 10;
// bram[7379] = 16;
// bram[7380] = 23;
// bram[7381] = 31;
// bram[7382] = 40;
// bram[7383] = 50;
// bram[7384] = 60;
// bram[7385] = 72;
// bram[7386] = 84;
// bram[7387] = 97;
// bram[7388] = 109;
// bram[7389] = 122;
// bram[7390] = 135;
// bram[7391] = 148;
// bram[7392] = 161;
// bram[7393] = 174;
// bram[7394] = 185;
// bram[7395] = 197;
// bram[7396] = 207;
// bram[7397] = 217;
// bram[7398] = 225;
// bram[7399] = 233;
// bram[7400] = 240;
// bram[7401] = 245;
// bram[7402] = 249;
// bram[7403] = 252;
// bram[7404] = 253;
// bram[7405] = 253;
// bram[7406] = 252;
// bram[7407] = 250;
// bram[7408] = 246;
// bram[7409] = 241;
// bram[7410] = 234;
// bram[7411] = 227;
// bram[7412] = 218;
// bram[7413] = 209;
// bram[7414] = 198;
// bram[7415] = 187;
// bram[7416] = 175;
// bram[7417] = 163;
// bram[7418] = 150;
// bram[7419] = 138;
// bram[7420] = 125;
// bram[7421] = 111;
// bram[7422] = 99;
// bram[7423] = 86;
// bram[7424] = 74;
// bram[7425] = 62;
// bram[7426] = 51;
// bram[7427] = 41;
// bram[7428] = 32;
// bram[7429] = 24;
// bram[7430] = 17;
// bram[7431] = 11;
// bram[7432] = 6;
// bram[7433] = 2;
// bram[7434] = 0;
// bram[7435] = 0;
// bram[7436] = 0;
// bram[7437] = 2;
// bram[7438] = 5;
// bram[7439] = 10;
// bram[7440] = 15;
// bram[7441] = 22;
// bram[7442] = 30;
// bram[7443] = 39;
// bram[7444] = 49;
// bram[7445] = 60;
// bram[7446] = 71;
// bram[7447] = 83;
// bram[7448] = 96;
// bram[7449] = 109;
// bram[7450] = 122;
// bram[7451] = 135;
// bram[7452] = 148;
// bram[7453] = 160;
// bram[7454] = 173;
// bram[7455] = 185;
// bram[7456] = 196;
// bram[7457] = 206;
// bram[7458] = 216;
// bram[7459] = 225;
// bram[7460] = 233;
// bram[7461] = 239;
// bram[7462] = 245;
// bram[7463] = 249;
// bram[7464] = 252;
// bram[7465] = 253;
// bram[7466] = 253;
// bram[7467] = 252;
// bram[7468] = 250;
// bram[7469] = 246;
// bram[7470] = 241;
// bram[7471] = 235;
// bram[7472] = 227;
// bram[7473] = 219;
// bram[7474] = 209;
// bram[7475] = 199;
// bram[7476] = 188;
// bram[7477] = 176;
// bram[7478] = 164;
// bram[7479] = 151;
// bram[7480] = 138;
// bram[7481] = 125;
// bram[7482] = 112;
// bram[7483] = 99;
// bram[7484] = 87;
// bram[7485] = 75;
// bram[7486] = 63;
// bram[7487] = 52;
// bram[7488] = 42;
// bram[7489] = 33;
// bram[7490] = 24;
// bram[7491] = 17;
// bram[7492] = 11;
// bram[7493] = 6;
// bram[7494] = 3;
// bram[7495] = 0;
// bram[7496] = 0;
// bram[7497] = 0;
// bram[7498] = 2;
// bram[7499] = 5;
// bram[7500] = 9;
// bram[7501] = 15;
// bram[7502] = 22;
// bram[7503] = 29;
// bram[7504] = 38;
// bram[7505] = 48;
// bram[7506] = 59;
// bram[7507] = 70;
// bram[7508] = 82;
// bram[7509] = 95;
// bram[7510] = 108;
// bram[7511] = 121;
// bram[7512] = 134;
// bram[7513] = 147;
// bram[7514] = 159;
// bram[7515] = 172;
// bram[7516] = 184;
// bram[7517] = 195;
// bram[7518] = 206;
// bram[7519] = 216;
// bram[7520] = 224;
// bram[7521] = 232;
// bram[7522] = 239;
// bram[7523] = 244;
// bram[7524] = 249;
// bram[7525] = 252;
// bram[7526] = 253;
// bram[7527] = 253;
// bram[7528] = 252;
// bram[7529] = 250;
// bram[7530] = 246;
// bram[7531] = 241;
// bram[7532] = 235;
// bram[7533] = 228;
// bram[7534] = 219;
// bram[7535] = 210;
// bram[7536] = 200;
// bram[7537] = 189;
// bram[7538] = 177;
// bram[7539] = 165;
// bram[7540] = 152;
// bram[7541] = 139;
// bram[7542] = 126;
// bram[7543] = 113;
// bram[7544] = 100;
// bram[7545] = 88;
// bram[7546] = 76;
// bram[7547] = 64;
// bram[7548] = 53;
// bram[7549] = 43;
// bram[7550] = 33;
// bram[7551] = 25;
// bram[7552] = 18;
// bram[7553] = 11;
// bram[7554] = 7;
// bram[7555] = 3;
// bram[7556] = 1;
// bram[7557] = 0;
// bram[7558] = 0;
// bram[7559] = 2;
// bram[7560] = 5;
// bram[7561] = 9;
// bram[7562] = 14;
// bram[7563] = 21;
// bram[7564] = 29;
// bram[7565] = 38;
// bram[7566] = 48;
// bram[7567] = 58;
// bram[7568] = 70;
// bram[7569] = 82;
// bram[7570] = 94;
// bram[7571] = 107;
// bram[7572] = 120;
// bram[7573] = 133;
// bram[7574] = 146;
// bram[7575] = 159;
// bram[7576] = 171;
// bram[7577] = 183;
// bram[7578] = 194;
// bram[7579] = 205;
// bram[7580] = 215;
// bram[7581] = 224;
// bram[7582] = 232;
// bram[7583] = 238;
// bram[7584] = 244;
// bram[7585] = 248;
// bram[7586] = 251;
// bram[7587] = 253;
// bram[7588] = 253;
// bram[7589] = 253;
// bram[7590] = 250;
// bram[7591] = 247;
// bram[7592] = 242;
// bram[7593] = 236;
// bram[7594] = 228;
// bram[7595] = 220;
// bram[7596] = 211;
// bram[7597] = 201;
// bram[7598] = 190;
// bram[7599] = 178;
// bram[7600] = 166;
// bram[7601] = 153;
// bram[7602] = 140;
// bram[7603] = 127;
// bram[7604] = 114;
// bram[7605] = 101;
// bram[7606] = 89;
// bram[7607] = 76;
// bram[7608] = 65;
// bram[7609] = 54;
// bram[7610] = 43;
// bram[7611] = 34;
// bram[7612] = 25;
// bram[7613] = 18;
// bram[7614] = 12;
// bram[7615] = 7;
// bram[7616] = 3;
// bram[7617] = 1;
// bram[7618] = 0;
// bram[7619] = 0;
// bram[7620] = 1;
// bram[7621] = 4;
// bram[7622] = 8;
// bram[7623] = 14;
// bram[7624] = 21;
// bram[7625] = 28;
// bram[7626] = 37;
// bram[7627] = 47;
// bram[7628] = 57;
// bram[7629] = 69;
// bram[7630] = 81;
// bram[7631] = 93;
// bram[7632] = 106;
// bram[7633] = 119;
// bram[7634] = 132;
// bram[7635] = 145;
// bram[7636] = 158;
// bram[7637] = 170;
// bram[7638] = 182;
// bram[7639] = 194;
// bram[7640] = 204;
// bram[7641] = 214;
// bram[7642] = 223;
// bram[7643] = 231;
// bram[7644] = 238;
// bram[7645] = 244;
// bram[7646] = 248;
// bram[7647] = 251;
// bram[7648] = 253;
// bram[7649] = 253;
// bram[7650] = 253;
// bram[7651] = 250;
// bram[7652] = 247;
// bram[7653] = 242;
// bram[7654] = 236;
// bram[7655] = 229;
// bram[7656] = 221;
// bram[7657] = 211;
// bram[7658] = 201;
// bram[7659] = 190;
// bram[7660] = 179;
// bram[7661] = 167;
// bram[7662] = 154;
// bram[7663] = 141;
// bram[7664] = 128;
// bram[7665] = 115;
// bram[7666] = 102;
// bram[7667] = 89;
// bram[7668] = 77;
// bram[7669] = 65;
// bram[7670] = 54;
// bram[7671] = 44;
// bram[7672] = 34;
// bram[7673] = 26;
// bram[7674] = 19;
// bram[7675] = 12;
// bram[7676] = 7;
// bram[7677] = 3;
// bram[7678] = 1;
// bram[7679] = 0;
// bram[7680] = 0;
// bram[7681] = 1;
// bram[7682] = 4;
// bram[7683] = 8;
// bram[7684] = 14;
// bram[7685] = 20;
// bram[7686] = 28;
// bram[7687] = 36;
// bram[7688] = 46;
// bram[7689] = 57;
// bram[7690] = 68;
// bram[7691] = 80;
// bram[7692] = 92;
// bram[7693] = 105;
// bram[7694] = 118;
// bram[7695] = 131;
// bram[7696] = 144;
// bram[7697] = 157;
// bram[7698] = 169;
// bram[7699] = 181;
// bram[7700] = 193;
// bram[7701] = 204;
// bram[7702] = 214;
// bram[7703] = 223;
// bram[7704] = 231;
// bram[7705] = 238;
// bram[7706] = 243;
// bram[7707] = 248;
// bram[7708] = 251;
// bram[7709] = 253;
// bram[7710] = 253;
// bram[7711] = 253;
// bram[7712] = 251;
// bram[7713] = 247;
// bram[7714] = 242;
// bram[7715] = 237;
// bram[7716] = 229;
// bram[7717] = 221;
// bram[7718] = 212;
// bram[7719] = 202;
// bram[7720] = 191;
// bram[7721] = 180;
// bram[7722] = 167;
// bram[7723] = 155;
// bram[7724] = 142;
// bram[7725] = 129;
// bram[7726] = 116;
// bram[7727] = 103;
// bram[7728] = 90;
// bram[7729] = 78;
// bram[7730] = 66;
// bram[7731] = 55;
// bram[7732] = 45;
// bram[7733] = 35;
// bram[7734] = 27;
// bram[7735] = 19;
// bram[7736] = 13;
// bram[7737] = 7;
// bram[7738] = 4;
// bram[7739] = 1;
// bram[7740] = 0;
// bram[7741] = 0;
// bram[7742] = 1;
// bram[7743] = 4;
// bram[7744] = 8;
// bram[7745] = 13;
// bram[7746] = 20;
// bram[7747] = 27;
// bram[7748] = 36;
// bram[7749] = 45;
// bram[7750] = 56;
// bram[7751] = 67;
// bram[7752] = 79;
// bram[7753] = 91;
// bram[7754] = 104;
// bram[7755] = 117;
// bram[7756] = 130;
// bram[7757] = 143;
// bram[7758] = 156;
// bram[7759] = 168;
// bram[7760] = 181;
// bram[7761] = 192;
// bram[7762] = 203;
// bram[7763] = 213;
// bram[7764] = 222;
// bram[7765] = 230;
// bram[7766] = 237;
// bram[7767] = 243;
// bram[7768] = 248;
// bram[7769] = 251;
// bram[7770] = 253;
// bram[7771] = 253;
// bram[7772] = 253;
// bram[7773] = 251;
// bram[7774] = 247;
// bram[7775] = 243;
// bram[7776] = 237;
// bram[7777] = 230;
// bram[7778] = 222;
// bram[7779] = 213;
// bram[7780] = 203;
// bram[7781] = 192;
// bram[7782] = 180;
// bram[7783] = 168;
// bram[7784] = 156;
// bram[7785] = 143;
// bram[7786] = 130;
// bram[7787] = 117;
// bram[7788] = 104;
// bram[7789] = 91;
// bram[7790] = 79;
// bram[7791] = 67;
// bram[7792] = 56;
// bram[7793] = 45;
// bram[7794] = 36;
// bram[7795] = 27;
// bram[7796] = 19;
// bram[7797] = 13;
// bram[7798] = 8;
// bram[7799] = 4;
// bram[7800] = 1;
// bram[7801] = 0;
// bram[7802] = 0;
// bram[7803] = 1;
// bram[7804] = 4;
// bram[7805] = 8;
// bram[7806] = 13;
// bram[7807] = 19;
// bram[7808] = 27;
// bram[7809] = 35;
// bram[7810] = 45;
// bram[7811] = 55;
// bram[7812] = 66;
// bram[7813] = 78;
// bram[7814] = 90;
// bram[7815] = 103;
// bram[7816] = 116;
// bram[7817] = 129;
// bram[7818] = 142;
// bram[7819] = 155;
// bram[7820] = 168;
// bram[7821] = 180;
// bram[7822] = 191;
// bram[7823] = 202;
// bram[7824] = 212;
// bram[7825] = 221;
// bram[7826] = 230;
// bram[7827] = 237;
// bram[7828] = 243;
// bram[7829] = 247;
// bram[7830] = 251;
// bram[7831] = 253;
// bram[7832] = 253;
// bram[7833] = 253;
// bram[7834] = 251;
// bram[7835] = 248;
// bram[7836] = 243;
// bram[7837] = 237;
// bram[7838] = 231;
// bram[7839] = 222;
// bram[7840] = 213;
// bram[7841] = 203;
// bram[7842] = 193;
// bram[7843] = 181;
// bram[7844] = 169;
// bram[7845] = 157;
// bram[7846] = 144;
// bram[7847] = 131;
// bram[7848] = 118;
// bram[7849] = 105;
// bram[7850] = 92;
// bram[7851] = 80;
// bram[7852] = 68;
// bram[7853] = 57;
// bram[7854] = 46;
// bram[7855] = 36;
// bram[7856] = 28;
// bram[7857] = 20;
// bram[7858] = 13;
// bram[7859] = 8;
// bram[7860] = 4;
// bram[7861] = 1;
// bram[7862] = 0;
// bram[7863] = 0;
// bram[7864] = 1;
// bram[7865] = 3;
// bram[7866] = 7;
// bram[7867] = 12;
// bram[7868] = 19;
// bram[7869] = 26;
// bram[7870] = 35;
// bram[7871] = 44;
// bram[7872] = 54;
// bram[7873] = 66;
// bram[7874] = 77;
// bram[7875] = 90;
// bram[7876] = 102;
// bram[7877] = 115;
// bram[7878] = 128;
// bram[7879] = 141;
// bram[7880] = 154;
// bram[7881] = 167;
// bram[7882] = 179;
// bram[7883] = 191;
// bram[7884] = 201;
// bram[7885] = 212;
// bram[7886] = 221;
// bram[7887] = 229;
// bram[7888] = 236;
// bram[7889] = 242;
// bram[7890] = 247;
// bram[7891] = 250;
// bram[7892] = 253;
// bram[7893] = 253;
// bram[7894] = 253;
// bram[7895] = 251;
// bram[7896] = 248;
// bram[7897] = 244;
// bram[7898] = 238;
// bram[7899] = 231;
// bram[7900] = 223;
// bram[7901] = 214;
// bram[7902] = 204;
// bram[7903] = 193;
// bram[7904] = 182;
// bram[7905] = 170;
// bram[7906] = 158;
// bram[7907] = 145;
// bram[7908] = 132;
// bram[7909] = 119;
// bram[7910] = 106;
// bram[7911] = 93;
// bram[7912] = 80;
// bram[7913] = 69;
// bram[7914] = 57;
// bram[7915] = 47;
// bram[7916] = 37;
// bram[7917] = 28;
// bram[7918] = 20;
// bram[7919] = 14;
// bram[7920] = 8;
// bram[7921] = 4;
// bram[7922] = 1;
// bram[7923] = 0;
// bram[7924] = 0;
// bram[7925] = 1;
// bram[7926] = 3;
// bram[7927] = 7;
// bram[7928] = 12;
// bram[7929] = 18;
// bram[7930] = 26;
// bram[7931] = 34;
// bram[7932] = 43;
// bram[7933] = 54;
// bram[7934] = 65;
// bram[7935] = 77;
// bram[7936] = 89;
// bram[7937] = 101;
// bram[7938] = 114;
// bram[7939] = 127;
// bram[7940] = 140;
// bram[7941] = 153;
// bram[7942] = 166;
// bram[7943] = 178;
// bram[7944] = 190;
// bram[7945] = 201;
// bram[7946] = 211;
// bram[7947] = 220;
// bram[7948] = 229;
// bram[7949] = 236;
// bram[7950] = 242;
// bram[7951] = 247;
// bram[7952] = 250;
// bram[7953] = 253;
// bram[7954] = 253;
// bram[7955] = 253;
// bram[7956] = 251;
// bram[7957] = 248;
// bram[7958] = 244;
// bram[7959] = 238;
// bram[7960] = 232;
// bram[7961] = 224;
// bram[7962] = 215;
// bram[7963] = 205;
// bram[7964] = 194;
// bram[7965] = 183;
// bram[7966] = 171;
// bram[7967] = 158;
// bram[7968] = 146;
// bram[7969] = 133;
// bram[7970] = 120;
// bram[7971] = 107;
// bram[7972] = 94;
// bram[7973] = 81;
// bram[7974] = 69;
// bram[7975] = 58;
// bram[7976] = 47;
// bram[7977] = 38;
// bram[7978] = 29;
// bram[7979] = 21;
// bram[7980] = 14;
// bram[7981] = 9;
// bram[7982] = 4;
// bram[7983] = 2;
// bram[7984] = 0;
// bram[7985] = 0;
// bram[7986] = 1;
// bram[7987] = 3;
// bram[7988] = 7;
// bram[7989] = 12;
// bram[7990] = 18;
// bram[7991] = 25;
// bram[7992] = 33;
// bram[7993] = 43;
// bram[7994] = 53;
// bram[7995] = 64;
// bram[7996] = 76;
// bram[7997] = 88;
// bram[7998] = 101;
// bram[7999] = 113;
// bram[8000] = 127;
// bram[8001] = 141;
// bram[8002] = 156;
// bram[8003] = 170;
// bram[8004] = 183;
// bram[8005] = 196;
// bram[8006] = 208;
// bram[8007] = 218;
// bram[8008] = 228;
// bram[8009] = 236;
// bram[8010] = 243;
// bram[8011] = 248;
// bram[8012] = 251;
// bram[8013] = 253;
// bram[8014] = 253;
// bram[8015] = 252;
// bram[8016] = 249;
// bram[8017] = 244;
// bram[8018] = 238;
// bram[8019] = 230;
// bram[8020] = 220;
// bram[8021] = 210;
// bram[8022] = 198;
// bram[8023] = 186;
// bram[8024] = 173;
// bram[8025] = 159;
// bram[8026] = 144;
// bram[8027] = 130;
// bram[8028] = 115;
// bram[8029] = 100;
// bram[8030] = 86;
// bram[8031] = 73;
// bram[8032] = 60;
// bram[8033] = 48;
// bram[8034] = 37;
// bram[8035] = 27;
// bram[8036] = 19;
// bram[8037] = 12;
// bram[8038] = 6;
// bram[8039] = 2;
// bram[8040] = 0;
// bram[8041] = 0;
// bram[8042] = 1;
// bram[8043] = 4;
// bram[8044] = 8;
// bram[8045] = 14;
// bram[8046] = 22;
// bram[8047] = 31;
// bram[8048] = 41;
// bram[8049] = 52;
// bram[8050] = 64;
// bram[8051] = 78;
// bram[8052] = 91;
// bram[8053] = 106;
// bram[8054] = 120;
// bram[8055] = 135;
// bram[8056] = 150;
// bram[8057] = 164;
// bram[8058] = 177;
// bram[8059] = 191;
// bram[8060] = 203;
// bram[8061] = 214;
// bram[8062] = 224;
// bram[8063] = 233;
// bram[8064] = 240;
// bram[8065] = 246;
// bram[8066] = 250;
// bram[8067] = 253;
// bram[8068] = 253;
// bram[8069] = 253;
// bram[8070] = 250;
// bram[8071] = 246;
// bram[8072] = 240;
// bram[8073] = 233;
// bram[8074] = 224;
// bram[8075] = 215;
// bram[8076] = 203;
// bram[8077] = 191;
// bram[8078] = 178;
// bram[8079] = 165;
// bram[8080] = 150;
// bram[8081] = 136;
// bram[8082] = 121;
// bram[8083] = 107;
// bram[8084] = 92;
// bram[8085] = 78;
// bram[8086] = 65;
// bram[8087] = 53;
// bram[8088] = 41;
// bram[8089] = 31;
// bram[8090] = 22;
// bram[8091] = 14;
// bram[8092] = 8;
// bram[8093] = 4;
// bram[8094] = 1;
// bram[8095] = 0;
// bram[8096] = 0;
// bram[8097] = 2;
// bram[8098] = 6;
// bram[8099] = 11;
// bram[8100] = 18;
// bram[8101] = 27;
// bram[8102] = 36;
// bram[8103] = 47;
// bram[8104] = 59;
// bram[8105] = 72;
// bram[8106] = 86;
// bram[8107] = 100;
// bram[8108] = 114;
// bram[8109] = 129;
// bram[8110] = 143;
// bram[8111] = 158;
// bram[8112] = 172;
// bram[8113] = 185;
// bram[8114] = 198;
// bram[8115] = 209;
// bram[8116] = 220;
// bram[8117] = 229;
// bram[8118] = 237;
// bram[8119] = 244;
// bram[8120] = 248;
// bram[8121] = 252;
// bram[8122] = 253;
// bram[8123] = 253;
// bram[8124] = 251;
// bram[8125] = 248;
// bram[8126] = 243;
// bram[8127] = 236;
// bram[8128] = 228;
// bram[8129] = 219;
// bram[8130] = 208;
// bram[8131] = 196;
// bram[8132] = 184;
// bram[8133] = 170;
// bram[8134] = 156;
// bram[8135] = 142;
// bram[8136] = 127;
// bram[8137] = 113;
// bram[8138] = 98;
// bram[8139] = 84;
// bram[8140] = 71;
// bram[8141] = 58;
// bram[8142] = 46;
// bram[8143] = 35;
// bram[8144] = 26;
// bram[8145] = 17;
// bram[8146] = 11;
// bram[8147] = 5;
// bram[8148] = 2;
// bram[8149] = 0;
// bram[8150] = 0;
// bram[8151] = 1;
// bram[8152] = 4;
// bram[8153] = 9;
// bram[8154] = 15;
// bram[8155] = 23;
// bram[8156] = 32;
// bram[8157] = 42;
// bram[8158] = 54;
// bram[8159] = 66;
// bram[8160] = 80;
// bram[8161] = 94;
// bram[8162] = 108;
// bram[8163] = 123;
// bram[8164] = 137;
// bram[8165] = 152;
// bram[8166] = 166;
// bram[8167] = 180;
// bram[8168] = 193;
// bram[8169] = 205;
// bram[8170] = 216;
// bram[8171] = 225;
// bram[8172] = 234;
// bram[8173] = 241;
// bram[8174] = 247;
// bram[8175] = 251;
// bram[8176] = 253;
// bram[8177] = 253;
// bram[8178] = 252;
// bram[8179] = 250;
// bram[8180] = 245;
// bram[8181] = 239;
// bram[8182] = 232;
// bram[8183] = 223;
// bram[8184] = 213;
// bram[8185] = 202;
// bram[8186] = 189;
// bram[8187] = 176;
// bram[8188] = 162;
// bram[8189] = 148;
// bram[8190] = 133;
// bram[8191] = 119;
// bram[8192] = 104;
// bram[8193] = 90;
// bram[8194] = 76;
// bram[8195] = 63;
// bram[8196] = 51;
// bram[8197] = 40;
// bram[8198] = 30;
// bram[8199] = 21;
// bram[8200] = 13;
// bram[8201] = 7;
// bram[8202] = 3;
// bram[8203] = 0;
// bram[8204] = 0;
// bram[8205] = 0;
// bram[8206] = 3;
// bram[8207] = 7;
// bram[8208] = 12;
// bram[8209] = 19;
// bram[8210] = 28;
// bram[8211] = 38;
// bram[8212] = 49;
// bram[8213] = 61;
// bram[8214] = 74;
// bram[8215] = 88;
// bram[8216] = 102;
// bram[8217] = 116;
// bram[8218] = 131;
// bram[8219] = 146;
// bram[8220] = 160;
// bram[8221] = 174;
// bram[8222] = 187;
// bram[8223] = 200;
// bram[8224] = 211;
// bram[8225] = 221;
// bram[8226] = 231;
// bram[8227] = 238;
// bram[8228] = 244;
// bram[8229] = 249;
// bram[8230] = 252;
// bram[8231] = 253;
// bram[8232] = 253;
// bram[8233] = 251;
// bram[8234] = 247;
// bram[8235] = 242;
// bram[8236] = 235;
// bram[8237] = 227;
// bram[8238] = 217;
// bram[8239] = 206;
// bram[8240] = 195;
// bram[8241] = 182;
// bram[8242] = 168;
// bram[8243] = 154;
// bram[8244] = 140;
// bram[8245] = 125;
// bram[8246] = 110;
// bram[8247] = 96;
// bram[8248] = 82;
// bram[8249] = 69;
// bram[8250] = 56;
// bram[8251] = 44;
// bram[8252] = 34;
// bram[8253] = 24;
// bram[8254] = 16;
// bram[8255] = 10;
// bram[8256] = 5;
// bram[8257] = 1;
// bram[8258] = 0;
// bram[8259] = 0;
// bram[8260] = 1;
// bram[8261] = 5;
// bram[8262] = 10;
// bram[8263] = 16;
// bram[8264] = 24;
// bram[8265] = 34;
// bram[8266] = 44;
// bram[8267] = 56;
// bram[8268] = 68;
// bram[8269] = 82;
// bram[8270] = 96;
// bram[8271] = 110;
// bram[8272] = 125;
// bram[8273] = 140;
// bram[8274] = 154;
// bram[8275] = 168;
// bram[8276] = 182;
// bram[8277] = 194;
// bram[8278] = 206;
// bram[8279] = 217;
// bram[8280] = 227;
// bram[8281] = 235;
// bram[8282] = 242;
// bram[8283] = 247;
// bram[8284] = 251;
// bram[8285] = 253;
// bram[8286] = 253;
// bram[8287] = 252;
// bram[8288] = 249;
// bram[8289] = 244;
// bram[8290] = 238;
// bram[8291] = 231;
// bram[8292] = 221;
// bram[8293] = 211;
// bram[8294] = 200;
// bram[8295] = 187;
// bram[8296] = 174;
// bram[8297] = 160;
// bram[8298] = 146;
// bram[8299] = 131;
// bram[8300] = 117;
// bram[8301] = 102;
// bram[8302] = 88;
// bram[8303] = 74;
// bram[8304] = 61;
// bram[8305] = 49;
// bram[8306] = 38;
// bram[8307] = 28;
// bram[8308] = 19;
// bram[8309] = 12;
// bram[8310] = 7;
// bram[8311] = 3;
// bram[8312] = 0;
// bram[8313] = 0;
// bram[8314] = 0;
// bram[8315] = 3;
// bram[8316] = 7;
// bram[8317] = 13;
// bram[8318] = 21;
// bram[8319] = 29;
// bram[8320] = 40;
// bram[8321] = 51;
// bram[8322] = 63;
// bram[8323] = 76;
// bram[8324] = 90;
// bram[8325] = 104;
// bram[8326] = 119;
// bram[8327] = 133;
// bram[8328] = 148;
// bram[8329] = 162;
// bram[8330] = 176;
// bram[8331] = 189;
// bram[8332] = 201;
// bram[8333] = 213;
// bram[8334] = 223;
// bram[8335] = 232;
// bram[8336] = 239;
// bram[8337] = 245;
// bram[8338] = 250;
// bram[8339] = 252;
// bram[8340] = 253;
// bram[8341] = 253;
// bram[8342] = 251;
// bram[8343] = 247;
// bram[8344] = 241;
// bram[8345] = 234;
// bram[8346] = 225;
// bram[8347] = 216;
// bram[8348] = 205;
// bram[8349] = 193;
// bram[8350] = 180;
// bram[8351] = 166;
// bram[8352] = 152;
// bram[8353] = 137;
// bram[8354] = 123;
// bram[8355] = 108;
// bram[8356] = 94;
// bram[8357] = 80;
// bram[8358] = 67;
// bram[8359] = 54;
// bram[8360] = 43;
// bram[8361] = 32;
// bram[8362] = 23;
// bram[8363] = 15;
// bram[8364] = 9;
// bram[8365] = 4;
// bram[8366] = 1;
// bram[8367] = 0;
// bram[8368] = 0;
// bram[8369] = 2;
// bram[8370] = 5;
// bram[8371] = 11;
// bram[8372] = 17;
// bram[8373] = 26;
// bram[8374] = 35;
// bram[8375] = 46;
// bram[8376] = 58;
// bram[8377] = 71;
// bram[8378] = 84;
// bram[8379] = 98;
// bram[8380] = 113;
// bram[8381] = 127;
// bram[8382] = 142;
// bram[8383] = 156;
// bram[8384] = 170;
// bram[8385] = 184;
// bram[8386] = 196;
// bram[8387] = 208;
// bram[8388] = 219;
// bram[8389] = 228;
// bram[8390] = 236;
// bram[8391] = 243;
// bram[8392] = 248;
// bram[8393] = 251;
// bram[8394] = 253;
// bram[8395] = 253;
// bram[8396] = 252;
// bram[8397] = 248;
// bram[8398] = 244;
// bram[8399] = 237;
// bram[8400] = 229;
// bram[8401] = 220;
// bram[8402] = 209;
// bram[8403] = 198;
// bram[8404] = 185;
// bram[8405] = 172;
// bram[8406] = 158;
// bram[8407] = 144;
// bram[8408] = 129;
// bram[8409] = 114;
// bram[8410] = 100;
// bram[8411] = 86;
// bram[8412] = 72;
// bram[8413] = 59;
// bram[8414] = 47;
// bram[8415] = 36;
// bram[8416] = 27;
// bram[8417] = 18;
// bram[8418] = 11;
// bram[8419] = 6;
// bram[8420] = 2;
// bram[8421] = 0;
// bram[8422] = 0;
// bram[8423] = 1;
// bram[8424] = 4;
// bram[8425] = 8;
// bram[8426] = 14;
// bram[8427] = 22;
// bram[8428] = 31;
// bram[8429] = 41;
// bram[8430] = 53;
// bram[8431] = 65;
// bram[8432] = 78;
// bram[8433] = 92;
// bram[8434] = 106;
// bram[8435] = 121;
// bram[8436] = 136;
// bram[8437] = 150;
// bram[8438] = 164;
// bram[8439] = 178;
// bram[8440] = 191;
// bram[8441] = 203;
// bram[8442] = 214;
// bram[8443] = 224;
// bram[8444] = 233;
// bram[8445] = 240;
// bram[8446] = 246;
// bram[8447] = 250;
// bram[8448] = 253;
// bram[8449] = 253;
// bram[8450] = 253;
// bram[8451] = 250;
// bram[8452] = 246;
// bram[8453] = 240;
// bram[8454] = 233;
// bram[8455] = 224;
// bram[8456] = 214;
// bram[8457] = 203;
// bram[8458] = 191;
// bram[8459] = 178;
// bram[8460] = 164;
// bram[8461] = 150;
// bram[8462] = 135;
// bram[8463] = 120;
// bram[8464] = 106;
// bram[8465] = 92;
// bram[8466] = 78;
// bram[8467] = 65;
// bram[8468] = 52;
// bram[8469] = 41;
// bram[8470] = 31;
// bram[8471] = 22;
// bram[8472] = 14;
// bram[8473] = 8;
// bram[8474] = 4;
// bram[8475] = 1;
// bram[8476] = 0;
// bram[8477] = 0;
// bram[8478] = 2;
// bram[8479] = 6;
// bram[8480] = 12;
// bram[8481] = 19;
// bram[8482] = 27;
// bram[8483] = 37;
// bram[8484] = 48;
// bram[8485] = 60;
// bram[8486] = 73;
// bram[8487] = 86;
// bram[8488] = 100;
// bram[8489] = 115;
// bram[8490] = 129;
// bram[8491] = 144;
// bram[8492] = 158;
// bram[8493] = 172;
// bram[8494] = 186;
// bram[8495] = 198;
// bram[8496] = 210;
// bram[8497] = 220;
// bram[8498] = 230;
// bram[8499] = 237;
// bram[8500] = 244;
// bram[8501] = 249;
// bram[8502] = 252;
// bram[8503] = 253;
// bram[8504] = 253;
// bram[8505] = 251;
// bram[8506] = 248;
// bram[8507] = 243;
// bram[8508] = 236;
// bram[8509] = 228;
// bram[8510] = 218;
// bram[8511] = 208;
// bram[8512] = 196;
// bram[8513] = 183;
// bram[8514] = 170;
// bram[8515] = 156;
// bram[8516] = 141;
// bram[8517] = 127;
// bram[8518] = 112;
// bram[8519] = 98;
// bram[8520] = 83;
// bram[8521] = 70;
// bram[8522] = 57;
// bram[8523] = 45;
// bram[8524] = 35;
// bram[8525] = 25;
// bram[8526] = 17;
// bram[8527] = 10;
// bram[8528] = 5;
// bram[8529] = 2;
// bram[8530] = 0;
// bram[8531] = 0;
// bram[8532] = 1;
// bram[8533] = 4;
// bram[8534] = 9;
// bram[8535] = 15;
// bram[8536] = 23;
// bram[8537] = 32;
// bram[8538] = 43;
// bram[8539] = 55;
// bram[8540] = 67;
// bram[8541] = 80;
// bram[8542] = 94;
// bram[8543] = 109;
// bram[8544] = 123;
// bram[8545] = 138;
// bram[8546] = 152;
// bram[8547] = 167;
// bram[8548] = 180;
// bram[8549] = 193;
// bram[8550] = 205;
// bram[8551] = 216;
// bram[8552] = 226;
// bram[8553] = 234;
// bram[8554] = 241;
// bram[8555] = 247;
// bram[8556] = 251;
// bram[8557] = 253;
// bram[8558] = 253;
// bram[8559] = 252;
// bram[8560] = 250;
// bram[8561] = 245;
// bram[8562] = 239;
// bram[8563] = 231;
// bram[8564] = 223;
// bram[8565] = 212;
// bram[8566] = 201;
// bram[8567] = 189;
// bram[8568] = 175;
// bram[8569] = 162;
// bram[8570] = 147;
// bram[8571] = 133;
// bram[8572] = 118;
// bram[8573] = 104;
// bram[8574] = 89;
// bram[8575] = 76;
// bram[8576] = 63;
// bram[8577] = 50;
// bram[8578] = 39;
// bram[8579] = 29;
// bram[8580] = 20;
// bram[8581] = 13;
// bram[8582] = 7;
// bram[8583] = 3;
// bram[8584] = 0;
// bram[8585] = 0;
// bram[8586] = 0;
// bram[8587] = 3;
// bram[8588] = 7;
// bram[8589] = 13;
// bram[8590] = 20;
// bram[8591] = 28;
// bram[8592] = 38;
// bram[8593] = 50;
// bram[8594] = 62;
// bram[8595] = 75;
// bram[8596] = 88;
// bram[8597] = 103;
// bram[8598] = 117;
// bram[8599] = 132;
// bram[8600] = 146;
// bram[8601] = 161;
// bram[8602] = 175;
// bram[8603] = 188;
// bram[8604] = 200;
// bram[8605] = 212;
// bram[8606] = 222;
// bram[8607] = 231;
// bram[8608] = 239;
// bram[8609] = 245;
// bram[8610] = 249;
// bram[8611] = 252;
// bram[8612] = 253;
// bram[8613] = 253;
// bram[8614] = 251;
// bram[8615] = 247;
// bram[8616] = 242;
// bram[8617] = 235;
// bram[8618] = 226;
// bram[8619] = 217;
// bram[8620] = 206;
// bram[8621] = 194;
// bram[8622] = 181;
// bram[8623] = 168;
// bram[8624] = 153;
// bram[8625] = 139;
// bram[8626] = 124;
// bram[8627] = 110;
// bram[8628] = 95;
// bram[8629] = 81;
// bram[8630] = 68;
// bram[8631] = 55;
// bram[8632] = 44;
// bram[8633] = 33;
// bram[8634] = 24;
// bram[8635] = 16;
// bram[8636] = 9;
// bram[8637] = 5;
// bram[8638] = 1;
// bram[8639] = 0;
// bram[8640] = 0;
// bram[8641] = 2;
// bram[8642] = 5;
// bram[8643] = 10;
// bram[8644] = 17;
// bram[8645] = 25;
// bram[8646] = 34;
// bram[8647] = 45;
// bram[8648] = 56;
// bram[8649] = 69;
// bram[8650] = 83;
// bram[8651] = 97;
// bram[8652] = 111;
// bram[8653] = 126;
// bram[8654] = 140;
// bram[8655] = 155;
// bram[8656] = 169;
// bram[8657] = 182;
// bram[8658] = 195;
// bram[8659] = 207;
// bram[8660] = 218;
// bram[8661] = 227;
// bram[8662] = 236;
// bram[8663] = 242;
// bram[8664] = 248;
// bram[8665] = 251;
// bram[8666] = 253;
// bram[8667] = 253;
// bram[8668] = 252;
// bram[8669] = 249;
// bram[8670] = 244;
// bram[8671] = 238;
// bram[8672] = 230;
// bram[8673] = 221;
// bram[8674] = 211;
// bram[8675] = 199;
// bram[8676] = 187;
// bram[8677] = 173;
// bram[8678] = 159;
// bram[8679] = 145;
// bram[8680] = 130;
// bram[8681] = 116;
// bram[8682] = 101;
// bram[8683] = 87;
// bram[8684] = 74;
// bram[8685] = 61;
// bram[8686] = 49;
// bram[8687] = 37;
// bram[8688] = 28;
// bram[8689] = 19;
// bram[8690] = 12;
// bram[8691] = 6;
// bram[8692] = 2;
// bram[8693] = 0;
// bram[8694] = 0;
// bram[8695] = 1;
// bram[8696] = 3;
// bram[8697] = 8;
// bram[8698] = 14;
// bram[8699] = 21;
// bram[8700] = 30;
// bram[8701] = 40;
// bram[8702] = 51;
// bram[8703] = 64;
// bram[8704] = 77;
// bram[8705] = 91;
// bram[8706] = 105;
// bram[8707] = 119;
// bram[8708] = 134;
// bram[8709] = 149;
// bram[8710] = 163;
// bram[8711] = 177;
// bram[8712] = 190;
// bram[8713] = 202;
// bram[8714] = 213;
// bram[8715] = 223;
// bram[8716] = 232;
// bram[8717] = 240;
// bram[8718] = 246;
// bram[8719] = 250;
// bram[8720] = 252;
// bram[8721] = 253;
// bram[8722] = 253;
// bram[8723] = 250;
// bram[8724] = 246;
// bram[8725] = 241;
// bram[8726] = 234;
// bram[8727] = 225;
// bram[8728] = 215;
// bram[8729] = 204;
// bram[8730] = 192;
// bram[8731] = 179;
// bram[8732] = 165;
// bram[8733] = 151;
// bram[8734] = 137;
// bram[8735] = 122;
// bram[8736] = 107;
// bram[8737] = 93;
// bram[8738] = 79;
// bram[8739] = 66;
// bram[8740] = 53;
// bram[8741] = 42;
// bram[8742] = 32;
// bram[8743] = 23;
// bram[8744] = 15;
// bram[8745] = 9;
// bram[8746] = 4;
// bram[8747] = 1;
// bram[8748] = 0;
// bram[8749] = 0;
// bram[8750] = 2;
// bram[8751] = 6;
// bram[8752] = 11;
// bram[8753] = 18;
// bram[8754] = 26;
// bram[8755] = 36;
// bram[8756] = 46;
// bram[8757] = 58;
// bram[8758] = 71;
// bram[8759] = 85;
// bram[8760] = 99;
// bram[8761] = 113;
// bram[8762] = 128;
// bram[8763] = 143;
// bram[8764] = 157;
// bram[8765] = 171;
// bram[8766] = 184;
// bram[8767] = 197;
// bram[8768] = 209;
// bram[8769] = 219;
// bram[8770] = 229;
// bram[8771] = 237;
// bram[8772] = 243;
// bram[8773] = 248;
// bram[8774] = 252;
// bram[8775] = 253;
// bram[8776] = 253;
// bram[8777] = 252;
// bram[8778] = 248;
// bram[8779] = 243;
// bram[8780] = 237;
// bram[8781] = 229;
// bram[8782] = 219;
// bram[8783] = 209;
// bram[8784] = 197;
// bram[8785] = 185;
// bram[8786] = 171;
// bram[8787] = 157;
// bram[8788] = 143;
// bram[8789] = 128;
// bram[8790] = 114;
// bram[8791] = 99;
// bram[8792] = 85;
// bram[8793] = 71;
// bram[8794] = 59;
// bram[8795] = 47;
// bram[8796] = 36;
// bram[8797] = 26;
// bram[8798] = 18;
// bram[8799] = 11;
// bram[8800] = 6;
// bram[8801] = 2;
// bram[8802] = 0;
// bram[8803] = 0;
// bram[8804] = 1;
// bram[8805] = 4;
// bram[8806] = 8;
// bram[8807] = 15;
// bram[8808] = 22;
// bram[8809] = 31;
// bram[8810] = 42;
// bram[8811] = 53;
// bram[8812] = 66;
// bram[8813] = 79;
// bram[8814] = 93;
// bram[8815] = 107;
// bram[8816] = 122;
// bram[8817] = 136;
// bram[8818] = 151;
// bram[8819] = 165;
// bram[8820] = 179;
// bram[8821] = 192;
// bram[8822] = 204;
// bram[8823] = 215;
// bram[8824] = 225;
// bram[8825] = 233;
// bram[8826] = 241;
// bram[8827] = 246;
// bram[8828] = 250;
// bram[8829] = 253;
// bram[8830] = 253;
// bram[8831] = 253;
// bram[8832] = 250;
// bram[8833] = 246;
// bram[8834] = 240;
// bram[8835] = 232;
// bram[8836] = 224;
// bram[8837] = 214;
// bram[8838] = 202;
// bram[8839] = 190;
// bram[8840] = 177;
// bram[8841] = 163;
// bram[8842] = 149;
// bram[8843] = 134;
// bram[8844] = 120;
// bram[8845] = 105;
// bram[8846] = 91;
// bram[8847] = 77;
// bram[8848] = 64;
// bram[8849] = 52;
// bram[8850] = 40;
// bram[8851] = 30;
// bram[8852] = 21;
// bram[8853] = 14;
// bram[8854] = 8;
// bram[8855] = 3;
// bram[8856] = 1;
// bram[8857] = 0;
// bram[8858] = 0;
// bram[8859] = 2;
// bram[8860] = 6;
// bram[8861] = 12;
// bram[8862] = 19;
// bram[8863] = 27;
// bram[8864] = 37;
// bram[8865] = 48;
// bram[8866] = 60;
// bram[8867] = 73;
// bram[8868] = 87;
// bram[8869] = 101;
// bram[8870] = 116;
// bram[8871] = 130;
// bram[8872] = 145;
// bram[8873] = 159;
// bram[8874] = 173;
// bram[8875] = 186;
// bram[8876] = 199;
// bram[8877] = 210;
// bram[8878] = 221;
// bram[8879] = 230;
// bram[8880] = 238;
// bram[8881] = 244;
// bram[8882] = 249;
// bram[8883] = 252;
// bram[8884] = 253;
// bram[8885] = 253;
// bram[8886] = 251;
// bram[8887] = 248;
// bram[8888] = 242;
// bram[8889] = 236;
// bram[8890] = 227;
// bram[8891] = 218;
// bram[8892] = 207;
// bram[8893] = 195;
// bram[8894] = 183;
// bram[8895] = 169;
// bram[8896] = 155;
// bram[8897] = 141;
// bram[8898] = 126;
// bram[8899] = 111;
// bram[8900] = 97;
// bram[8901] = 83;
// bram[8902] = 69;
// bram[8903] = 57;
// bram[8904] = 45;
// bram[8905] = 34;
// bram[8906] = 25;
// bram[8907] = 17;
// bram[8908] = 10;
// bram[8909] = 5;
// bram[8910] = 2;
// bram[8911] = 0;
// bram[8912] = 0;
// bram[8913] = 1;
// bram[8914] = 4;
// bram[8915] = 9;
// bram[8916] = 16;
// bram[8917] = 24;
// bram[8918] = 33;
// bram[8919] = 43;
// bram[8920] = 55;
// bram[8921] = 68;
// bram[8922] = 81;
// bram[8923] = 95;
// bram[8924] = 109;
// bram[8925] = 124;
// bram[8926] = 139;
// bram[8927] = 153;
// bram[8928] = 167;
// bram[8929] = 181;
// bram[8930] = 194;
// bram[8931] = 206;
// bram[8932] = 217;
// bram[8933] = 226;
// bram[8934] = 235;
// bram[8935] = 242;
// bram[8936] = 247;
// bram[8937] = 251;
// bram[8938] = 253;
// bram[8939] = 253;
// bram[8940] = 252;
// bram[8941] = 249;
// bram[8942] = 245;
// bram[8943] = 239;
// bram[8944] = 231;
// bram[8945] = 222;
// bram[8946] = 212;
// bram[8947] = 200;
// bram[8948] = 188;
// bram[8949] = 175;
// bram[8950] = 161;
// bram[8951] = 147;
// bram[8952] = 132;
// bram[8953] = 117;
// bram[8954] = 103;
// bram[8955] = 89;
// bram[8956] = 75;
// bram[8957] = 62;
// bram[8958] = 50;
// bram[8959] = 39;
// bram[8960] = 29;
// bram[8961] = 20;
// bram[8962] = 13;
// bram[8963] = 7;
// bram[8964] = 3;
// bram[8965] = 0;
// bram[8966] = 0;
// bram[8967] = 0;
// bram[8968] = 3;
// bram[8969] = 7;
// bram[8970] = 13;
// bram[8971] = 20;
// bram[8972] = 29;
// bram[8973] = 39;
// bram[8974] = 50;
// bram[8975] = 62;
// bram[8976] = 75;
// bram[8977] = 89;
// bram[8978] = 103;
// bram[8979] = 118;
// bram[8980] = 132;
// bram[8981] = 147;
// bram[8982] = 161;
// bram[8983] = 175;
// bram[8984] = 188;
// bram[8985] = 201;
// bram[8986] = 212;
// bram[8987] = 222;
// bram[8988] = 231;
// bram[8989] = 239;
// bram[8990] = 245;
// bram[8991] = 249;
// bram[8992] = 252;
// bram[8993] = 253;
// bram[8994] = 253;
// bram[8995] = 251;
// bram[8996] = 247;
// bram[8997] = 241;
// bram[8998] = 234;
// bram[8999] = 226;
// bram[9000] = 216;
// bram[9001] = 205;
// bram[9002] = 193;
// bram[9003] = 180;
// bram[9004] = 167;
// bram[9005] = 153;
// bram[9006] = 138;
// bram[9007] = 124;
// bram[9008] = 109;
// bram[9009] = 95;
// bram[9010] = 81;
// bram[9011] = 67;
// bram[9012] = 55;
// bram[9013] = 43;
// bram[9014] = 33;
// bram[9015] = 23;
// bram[9016] = 16;
// bram[9017] = 9;
// bram[9018] = 4;
// bram[9019] = 1;
// bram[9020] = 0;
// bram[9021] = 0;
// bram[9022] = 2;
// bram[9023] = 5;
// bram[9024] = 10;
// bram[9025] = 17;
// bram[9026] = 25;
// bram[9027] = 35;
// bram[9028] = 45;
// bram[9029] = 57;
// bram[9030] = 70;
// bram[9031] = 83;
// bram[9032] = 97;
// bram[9033] = 112;
// bram[9034] = 126;
// bram[9035] = 141;
// bram[9036] = 155;
// bram[9037] = 169;
// bram[9038] = 183;
// bram[9039] = 196;
// bram[9040] = 207;
// bram[9041] = 218;
// bram[9042] = 228;
// bram[9043] = 236;
// bram[9044] = 243;
// bram[9045] = 248;
// bram[9046] = 251;
// bram[9047] = 253;
// bram[9048] = 253;
// bram[9049] = 252;
// bram[9050] = 249;
// bram[9051] = 244;
// bram[9052] = 238;
// bram[9053] = 230;
// bram[9054] = 221;
// bram[9055] = 210;
// bram[9056] = 199;
// bram[9057] = 186;
// bram[9058] = 173;
// bram[9059] = 159;
// bram[9060] = 144;
// bram[9061] = 130;
// bram[9062] = 115;
// bram[9063] = 101;
// bram[9064] = 86;
// bram[9065] = 73;
// bram[9066] = 60;
// bram[9067] = 48;
// bram[9068] = 37;
// bram[9069] = 27;
// bram[9070] = 19;
// bram[9071] = 12;
// bram[9072] = 6;
// bram[9073] = 2;
// bram[9074] = 0;
// bram[9075] = 0;
// bram[9076] = 1;
// bram[9077] = 3;
// bram[9078] = 8;
// bram[9079] = 14;
// bram[9080] = 21;
// bram[9081] = 30;
// bram[9082] = 41;
// bram[9083] = 52;
// bram[9084] = 64;
// bram[9085] = 77;
// bram[9086] = 91;
// bram[9087] = 106;
// bram[9088] = 120;
// bram[9089] = 135;
// bram[9090] = 149;
// bram[9091] = 164;
// bram[9092] = 177;
// bram[9093] = 190;
// bram[9094] = 203;
// bram[9095] = 214;
// bram[9096] = 224;
// bram[9097] = 233;
// bram[9098] = 240;
// bram[9099] = 246;
// bram[9100] = 250;
// bram[9101] = 253;
// bram[9102] = 253;
// bram[9103] = 253;
// bram[9104] = 250;
// bram[9105] = 246;
// bram[9106] = 240;
// bram[9107] = 233;
// bram[9108] = 225;
// bram[9109] = 215;
// bram[9110] = 204;
// bram[9111] = 191;
// bram[9112] = 178;
// bram[9113] = 165;
// bram[9114] = 150;
// bram[9115] = 136;
// bram[9116] = 121;
// bram[9117] = 107;
// bram[9118] = 92;
// bram[9119] = 79;
// bram[9120] = 65;
// bram[9121] = 53;
// bram[9122] = 41;
// bram[9123] = 31;
// bram[9124] = 22;
// bram[9125] = 14;
// bram[9126] = 8;
// bram[9127] = 4;
// bram[9128] = 1;
// bram[9129] = 0;
// bram[9130] = 0;
// bram[9131] = 2;
// bram[9132] = 6;
// bram[9133] = 11;
// bram[9134] = 18;
// bram[9135] = 26;
// bram[9136] = 36;
// bram[9137] = 47;
// bram[9138] = 59;
// bram[9139] = 72;
// bram[9140] = 85;
// bram[9141] = 99;
// bram[9142] = 114;
// bram[9143] = 129;
// bram[9144] = 143;
// bram[9145] = 158;
// bram[9146] = 172;
// bram[9147] = 185;
// bram[9148] = 198;
// bram[9149] = 209;
// bram[9150] = 220;
// bram[9151] = 229;
// bram[9152] = 237;
// bram[9153] = 243;
// bram[9154] = 248;
// bram[9155] = 252;
// bram[9156] = 253;
// bram[9157] = 253;
// bram[9158] = 252;
// bram[9159] = 248;
// bram[9160] = 243;
// bram[9161] = 236;
// bram[9162] = 228;
// bram[9163] = 219;
// bram[9164] = 208;
// bram[9165] = 197;
// bram[9166] = 184;
// bram[9167] = 171;
// bram[9168] = 157;
// bram[9169] = 142;
// bram[9170] = 127;
// bram[9171] = 113;
// bram[9172] = 98;
// bram[9173] = 84;
// bram[9174] = 71;
// bram[9175] = 58;
// bram[9176] = 46;
// bram[9177] = 35;
// bram[9178] = 26;
// bram[9179] = 18;
// bram[9180] = 11;
// bram[9181] = 6;
// bram[9182] = 2;
// bram[9183] = 0;
// bram[9184] = 0;
// bram[9185] = 1;
// bram[9186] = 4;
// bram[9187] = 9;
// bram[9188] = 15;
// bram[9189] = 23;
// bram[9190] = 32;
// bram[9191] = 42;
// bram[9192] = 54;
// bram[9193] = 66;
// bram[9194] = 80;
// bram[9195] = 93;
// bram[9196] = 108;
// bram[9197] = 122;
// bram[9198] = 137;
// bram[9199] = 152;
// bram[9200] = 166;
// bram[9201] = 179;
// bram[9202] = 192;
// bram[9203] = 204;
// bram[9204] = 215;
// bram[9205] = 225;
// bram[9206] = 234;
// bram[9207] = 241;
// bram[9208] = 247;
// bram[9209] = 251;
// bram[9210] = 253;
// bram[9211] = 253;
// bram[9212] = 252;
// bram[9213] = 250;
// bram[9214] = 245;
// bram[9215] = 239;
// bram[9216] = 232;
// bram[9217] = 223;
// bram[9218] = 213;
// bram[9219] = 202;
// bram[9220] = 189;
// bram[9221] = 176;
// bram[9222] = 163;
// bram[9223] = 148;
// bram[9224] = 134;
// bram[9225] = 119;
// bram[9226] = 104;
// bram[9227] = 90;
// bram[9228] = 76;
// bram[9229] = 63;
// bram[9230] = 51;
// bram[9231] = 40;
// bram[9232] = 30;
// bram[9233] = 21;
// bram[9234] = 13;
// bram[9235] = 8;
// bram[9236] = 3;
// bram[9237] = 1;
// bram[9238] = 0;
// bram[9239] = 0;
// bram[9240] = 3;
// bram[9241] = 7;
// bram[9242] = 12;
// bram[9243] = 19;
// bram[9244] = 28;
// bram[9245] = 38;
// bram[9246] = 49;
// bram[9247] = 61;
// bram[9248] = 74;
// bram[9249] = 88;
// bram[9250] = 102;
// bram[9251] = 116;
// bram[9252] = 131;
// bram[9253] = 145;
// bram[9254] = 160;
// bram[9255] = 174;
// bram[9256] = 187;
// bram[9257] = 199;
// bram[9258] = 211;
// bram[9259] = 221;
// bram[9260] = 230;
// bram[9261] = 238;
// bram[9262] = 244;
// bram[9263] = 249;
// bram[9264] = 252;
// bram[9265] = 253;
// bram[9266] = 253;
// bram[9267] = 251;
// bram[9268] = 247;
// bram[9269] = 242;
// bram[9270] = 235;
// bram[9271] = 227;
// bram[9272] = 217;
// bram[9273] = 207;
// bram[9274] = 195;
// bram[9275] = 182;
// bram[9276] = 168;
// bram[9277] = 154;
// bram[9278] = 140;
// bram[9279] = 125;
// bram[9280] = 111;
// bram[9281] = 96;
// bram[9282] = 82;
// bram[9283] = 69;
// bram[9284] = 56;
// bram[9285] = 44;
// bram[9286] = 34;
// bram[9287] = 24;
// bram[9288] = 16;
// bram[9289] = 10;
// bram[9290] = 5;
// bram[9291] = 1;
// bram[9292] = 0;
// bram[9293] = 0;
// bram[9294] = 1;
// bram[9295] = 5;
// bram[9296] = 10;
// bram[9297] = 16;
// bram[9298] = 24;
// bram[9299] = 33;
// bram[9300] = 44;
// bram[9301] = 56;
// bram[9302] = 68;
// bram[9303] = 82;
// bram[9304] = 96;
// bram[9305] = 110;
// bram[9306] = 125;
// bram[9307] = 139;
// bram[9308] = 154;
// bram[9309] = 168;
// bram[9310] = 181;
// bram[9311] = 194;
// bram[9312] = 206;
// bram[9313] = 217;
// bram[9314] = 227;
// bram[9315] = 235;
// bram[9316] = 242;
// bram[9317] = 247;
// bram[9318] = 251;
// bram[9319] = 253;
// bram[9320] = 253;
// bram[9321] = 252;
// bram[9322] = 249;
// bram[9323] = 245;
// bram[9324] = 238;
// bram[9325] = 231;
// bram[9326] = 222;
// bram[9327] = 211;
// bram[9328] = 200;
// bram[9329] = 187;
// bram[9330] = 174;
// bram[9331] = 160;
// bram[9332] = 146;
// bram[9333] = 131;
// bram[9334] = 117;
// bram[9335] = 102;
// bram[9336] = 88;
// bram[9337] = 74;
// bram[9338] = 61;
// bram[9339] = 49;
// bram[9340] = 38;
// bram[9341] = 28;
// bram[9342] = 20;
// bram[9343] = 12;
// bram[9344] = 7;
// bram[9345] = 3;
// bram[9346] = 0;
// bram[9347] = 0;
// bram[9348] = 0;
// bram[9349] = 3;
// bram[9350] = 7;
// bram[9351] = 13;
// bram[9352] = 21;
// bram[9353] = 29;
// bram[9354] = 39;
// bram[9355] = 51;
// bram[9356] = 63;
// bram[9357] = 76;
// bram[9358] = 90;
// bram[9359] = 104;
// bram[9360] = 119;
// bram[9361] = 133;
// bram[9362] = 148;
// bram[9363] = 162;
// bram[9364] = 176;
// bram[9365] = 189;
// bram[9366] = 201;
// bram[9367] = 213;
// bram[9368] = 223;
// bram[9369] = 232;
// bram[9370] = 239;
// bram[9371] = 245;
// bram[9372] = 250;
// bram[9373] = 252;
// bram[9374] = 253;
// bram[9375] = 253;
// bram[9376] = 251;
// bram[9377] = 247;
// bram[9378] = 241;
// bram[9379] = 234;
// bram[9380] = 226;
// bram[9381] = 216;
// bram[9382] = 205;
// bram[9383] = 193;
// bram[9384] = 180;
// bram[9385] = 166;
// bram[9386] = 152;
// bram[9387] = 138;
// bram[9388] = 123;
// bram[9389] = 108;
// bram[9390] = 94;
// bram[9391] = 80;
// bram[9392] = 67;
// bram[9393] = 54;
// bram[9394] = 43;
// bram[9395] = 32;
// bram[9396] = 23;
// bram[9397] = 15;
// bram[9398] = 9;
// bram[9399] = 4;
// bram[9400] = 1;
// bram[9401] = 0;
// bram[9402] = 0;
// bram[9403] = 2;
// bram[9404] = 5;
// bram[9405] = 11;
// bram[9406] = 17;
// bram[9407] = 25;
// bram[9408] = 35;
// bram[9409] = 46;
// bram[9410] = 58;
// bram[9411] = 70;
// bram[9412] = 84;
// bram[9413] = 98;
// bram[9414] = 112;
// bram[9415] = 127;
// bram[9416] = 142;
// bram[9417] = 156;
// bram[9418] = 170;
// bram[9419] = 184;
// bram[9420] = 196;
// bram[9421] = 208;
// bram[9422] = 219;
// bram[9423] = 228;
// bram[9424] = 236;
// bram[9425] = 243;
// bram[9426] = 248;
// bram[9427] = 251;
// bram[9428] = 253;
// bram[9429] = 253;
// bram[9430] = 252;
// bram[9431] = 249;
// bram[9432] = 244;
// bram[9433] = 237;
// bram[9434] = 229;
// bram[9435] = 220;
// bram[9436] = 210;
// bram[9437] = 198;
// bram[9438] = 185;
// bram[9439] = 172;
// bram[9440] = 158;
// bram[9441] = 144;
// bram[9442] = 129;
// bram[9443] = 114;
// bram[9444] = 100;
// bram[9445] = 86;
// bram[9446] = 72;
// bram[9447] = 59;
// bram[9448] = 47;
// bram[9449] = 36;
// bram[9450] = 27;
// bram[9451] = 18;
// bram[9452] = 11;
// bram[9453] = 6;
// bram[9454] = 2;
// bram[9455] = 0;
// bram[9456] = 0;
// bram[9457] = 1;
// bram[9458] = 4;
// bram[9459] = 8;
// bram[9460] = 14;
// bram[9461] = 22;
// bram[9462] = 31;
// bram[9463] = 41;
// bram[9464] = 52;
// bram[9465] = 65;
// bram[9466] = 78;
// bram[9467] = 92;
// bram[9468] = 106;
// bram[9469] = 121;
// bram[9470] = 135;
// bram[9471] = 150;
// bram[9472] = 164;
// bram[9473] = 178;
// bram[9474] = 191;
// bram[9475] = 203;
// bram[9476] = 214;
// bram[9477] = 224;
// bram[9478] = 233;
// bram[9479] = 240;
// bram[9480] = 246;
// bram[9481] = 250;
// bram[9482] = 253;
// bram[9483] = 253;
// bram[9484] = 253;
// bram[9485] = 250;
// bram[9486] = 246;
// bram[9487] = 240;
// bram[9488] = 233;
// bram[9489] = 224;
// bram[9490] = 214;
// bram[9491] = 203;
// bram[9492] = 191;
// bram[9493] = 178;
// bram[9494] = 164;
// bram[9495] = 150;
// bram[9496] = 135;
// bram[9497] = 121;
// bram[9498] = 106;
// bram[9499] = 92;
// bram[9500] = 78;
// bram[9501] = 65;
// bram[9502] = 52;
// bram[9503] = 41;
// bram[9504] = 31;
// bram[9505] = 22;
// bram[9506] = 14;
// bram[9507] = 8;
// bram[9508] = 4;
// bram[9509] = 1;
// bram[9510] = 0;
// bram[9511] = 0;
// bram[9512] = 2;
// bram[9513] = 6;
// bram[9514] = 12;
// bram[9515] = 18;
// bram[9516] = 27;
// bram[9517] = 37;
// bram[9518] = 48;
// bram[9519] = 60;
// bram[9520] = 72;
// bram[9521] = 86;
// bram[9522] = 100;
// bram[9523] = 115;
// bram[9524] = 129;
// bram[9525] = 144;
// bram[9526] = 158;
// bram[9527] = 172;
// bram[9528] = 186;
// bram[9529] = 198;
// bram[9530] = 210;
// bram[9531] = 220;
// bram[9532] = 229;
// bram[9533] = 237;
// bram[9534] = 244;
// bram[9535] = 249;
// bram[9536] = 252;
// bram[9537] = 253;
// bram[9538] = 253;
// bram[9539] = 251;
// bram[9540] = 248;
// bram[9541] = 243;
// bram[9542] = 236;
// bram[9543] = 228;
// bram[9544] = 219;
// bram[9545] = 208;
// bram[9546] = 196;
// bram[9547] = 183;
// bram[9548] = 170;
// bram[9549] = 156;
// bram[9550] = 141;
// bram[9551] = 127;
// bram[9552] = 112;
// bram[9553] = 98;
// bram[9554] = 84;
// bram[9555] = 70;
// bram[9556] = 57;
// bram[9557] = 46;
// bram[9558] = 35;
// bram[9559] = 25;
// bram[9560] = 17;
// bram[9561] = 10;
// bram[9562] = 5;
// bram[9563] = 2;
// bram[9564] = 0;
// bram[9565] = 0;
// bram[9566] = 1;
// bram[9567] = 4;
// bram[9568] = 9;
// bram[9569] = 15;
// bram[9570] = 23;
// bram[9571] = 32;
// bram[9572] = 43;
// bram[9573] = 54;
// bram[9574] = 67;
// bram[9575] = 80;
// bram[9576] = 94;
// bram[9577] = 109;
// bram[9578] = 123;
// bram[9579] = 138;
// bram[9580] = 152;
// bram[9581] = 166;
// bram[9582] = 180;
// bram[9583] = 193;
// bram[9584] = 205;
// bram[9585] = 216;
// bram[9586] = 226;
// bram[9587] = 234;
// bram[9588] = 241;
// bram[9589] = 247;
// bram[9590] = 251;
// bram[9591] = 253;
// bram[9592] = 253;
// bram[9593] = 252;
// bram[9594] = 250;
// bram[9595] = 245;
// bram[9596] = 239;
// bram[9597] = 232;
// bram[9598] = 223;
// bram[9599] = 212;
// bram[9600] = 201;
// bram[9601] = 189;
// bram[9602] = 176;
// bram[9603] = 162;
// bram[9604] = 148;
// bram[9605] = 133;
// bram[9606] = 118;
// bram[9607] = 104;
// bram[9608] = 90;
// bram[9609] = 76;
// bram[9610] = 63;
// bram[9611] = 50;
// bram[9612] = 39;
// bram[9613] = 29;
// bram[9614] = 20;
// bram[9615] = 13;
// bram[9616] = 7;
// bram[9617] = 3;
// bram[9618] = 0;
// bram[9619] = 0;
// bram[9620] = 0;
// bram[9621] = 3;
// bram[9622] = 7;
// bram[9623] = 12;
// bram[9624] = 20;
// bram[9625] = 28;
// bram[9626] = 38;
// bram[9627] = 49;
// bram[9628] = 62;
// bram[9629] = 75;
// bram[9630] = 88;
// bram[9631] = 102;
// bram[9632] = 117;
// bram[9633] = 132;
// bram[9634] = 146;
// bram[9635] = 160;
// bram[9636] = 174;
// bram[9637] = 188;
// bram[9638] = 200;
// bram[9639] = 211;
// bram[9640] = 222;
// bram[9641] = 231;
// bram[9642] = 238;
// bram[9643] = 245;
// bram[9644] = 249;
// bram[9645] = 252;
// bram[9646] = 253;
// bram[9647] = 253;
// bram[9648] = 251;
// bram[9649] = 247;
// bram[9650] = 242;
// bram[9651] = 235;
// bram[9652] = 227;
// bram[9653] = 217;
// bram[9654] = 206;
// bram[9655] = 194;
// bram[9656] = 181;
// bram[9657] = 168;
// bram[9658] = 154;
// bram[9659] = 139;
// bram[9660] = 125;
// bram[9661] = 110;
// bram[9662] = 95;
// bram[9663] = 82;
// bram[9664] = 68;
// bram[9665] = 56;
// bram[9666] = 44;
// bram[9667] = 33;
// bram[9668] = 24;
// bram[9669] = 16;
// bram[9670] = 10;
// bram[9671] = 5;
// bram[9672] = 1;
// bram[9673] = 0;
// bram[9674] = 0;
// bram[9675] = 1;
// bram[9676] = 5;
// bram[9677] = 10;
// bram[9678] = 16;
// bram[9679] = 25;
// bram[9680] = 34;
// bram[9681] = 45;
// bram[9682] = 56;
// bram[9683] = 69;
// bram[9684] = 82;
// bram[9685] = 96;
// bram[9686] = 111;
// bram[9687] = 125;
// bram[9688] = 140;
// bram[9689] = 154;
// bram[9690] = 169;
// bram[9691] = 182;
// bram[9692] = 195;
// bram[9693] = 207;
// bram[9694] = 218;
// bram[9695] = 227;
// bram[9696] = 235;
// bram[9697] = 242;
// bram[9698] = 247;
// bram[9699] = 251;
// bram[9700] = 253;
// bram[9701] = 253;
// bram[9702] = 252;
// bram[9703] = 249;
// bram[9704] = 244;
// bram[9705] = 238;
// bram[9706] = 230;
// bram[9707] = 221;
// bram[9708] = 211;
// bram[9709] = 199;
// bram[9710] = 187;
// bram[9711] = 174;
// bram[9712] = 160;
// bram[9713] = 145;
// bram[9714] = 131;
// bram[9715] = 116;
// bram[9716] = 102;
// bram[9717] = 87;
// bram[9718] = 74;
// bram[9719] = 61;
// bram[9720] = 49;
// bram[9721] = 38;
// bram[9722] = 28;
// bram[9723] = 19;
// bram[9724] = 12;
// bram[9725] = 7;
// bram[9726] = 3;
// bram[9727] = 0;
// bram[9728] = 0;
// bram[9729] = 1;
// bram[9730] = 3;
// bram[9731] = 8;
// bram[9732] = 14;
// bram[9733] = 21;
// bram[9734] = 30;
// bram[9735] = 40;
// bram[9736] = 51;
// bram[9737] = 63;
// bram[9738] = 77;
// bram[9739] = 90;
// bram[9740] = 105;
// bram[9741] = 119;
// bram[9742] = 134;
// bram[9743] = 148;
// bram[9744] = 163;
// bram[9745] = 176;
// bram[9746] = 190;
// bram[9747] = 202;
// bram[9748] = 213;
// bram[9749] = 223;
// bram[9750] = 232;
// bram[9751] = 240;
// bram[9752] = 245;
// bram[9753] = 250;
// bram[9754] = 252;
// bram[9755] = 253;
// bram[9756] = 253;
// bram[9757] = 250;
// bram[9758] = 246;
// bram[9759] = 241;
// bram[9760] = 234;
// bram[9761] = 225;
// bram[9762] = 215;
// bram[9763] = 204;
// bram[9764] = 192;
// bram[9765] = 179;
// bram[9766] = 166;
// bram[9767] = 151;
// bram[9768] = 137;
// bram[9769] = 122;
// bram[9770] = 108;
// bram[9771] = 93;
// bram[9772] = 79;
// bram[9773] = 66;
// bram[9774] = 54;
// bram[9775] = 42;
// bram[9776] = 32;
// bram[9777] = 23;
// bram[9778] = 15;
// bram[9779] = 9;
// bram[9780] = 4;
// bram[9781] = 1;
// bram[9782] = 0;
// bram[9783] = 0;
// bram[9784] = 2;
// bram[9785] = 6;
// bram[9786] = 11;
// bram[9787] = 18;
// bram[9788] = 26;
// bram[9789] = 36;
// bram[9790] = 46;
// bram[9791] = 58;
// bram[9792] = 71;
// bram[9793] = 85;
// bram[9794] = 99;
// bram[9795] = 113;
// bram[9796] = 128;
// bram[9797] = 142;
// bram[9798] = 157;
// bram[9799] = 171;
// bram[9800] = 184;
// bram[9801] = 197;
// bram[9802] = 209;
// bram[9803] = 219;
// bram[9804] = 229;
// bram[9805] = 237;
// bram[9806] = 243;
// bram[9807] = 248;
// bram[9808] = 252;
// bram[9809] = 253;
// bram[9810] = 253;
// bram[9811] = 252;
// bram[9812] = 248;
// bram[9813] = 243;
// bram[9814] = 237;
// bram[9815] = 229;
// bram[9816] = 220;
// bram[9817] = 209;
// bram[9818] = 197;
// bram[9819] = 185;
// bram[9820] = 171;
// bram[9821] = 157;
// bram[9822] = 143;
// bram[9823] = 128;
// bram[9824] = 114;
// bram[9825] = 99;
// bram[9826] = 85;
// bram[9827] = 72;
// bram[9828] = 59;
// bram[9829] = 47;
// bram[9830] = 36;
// bram[9831] = 26;
// bram[9832] = 18;
// bram[9833] = 11;
// bram[9834] = 6;
// bram[9835] = 2;
// bram[9836] = 0;
// bram[9837] = 0;
// bram[9838] = 1;
// bram[9839] = 4;
// bram[9840] = 8;
// bram[9841] = 15;
// bram[9842] = 22;
// bram[9843] = 31;
// bram[9844] = 42;
// bram[9845] = 53;
// bram[9846] = 65;
// bram[9847] = 79;
// bram[9848] = 93;
// bram[9849] = 107;
// bram[9850] = 122;
// bram[9851] = 136;
// bram[9852] = 151;
// bram[9853] = 165;
// bram[9854] = 179;
// bram[9855] = 192;
// bram[9856] = 204;
// bram[9857] = 215;
// bram[9858] = 225;
// bram[9859] = 233;
// bram[9860] = 241;
// bram[9861] = 246;
// bram[9862] = 250;
// bram[9863] = 253;
// bram[9864] = 253;
// bram[9865] = 253;
// bram[9866] = 250;
// bram[9867] = 246;
// bram[9868] = 240;
// bram[9869] = 232;
// bram[9870] = 224;
// bram[9871] = 214;
// bram[9872] = 202;
// bram[9873] = 190;
// bram[9874] = 177;
// bram[9875] = 163;
// bram[9876] = 149;
// bram[9877] = 135;
// bram[9878] = 120;
// bram[9879] = 105;
// bram[9880] = 91;
// bram[9881] = 77;
// bram[9882] = 64;
// bram[9883] = 52;
// bram[9884] = 40;
// bram[9885] = 30;
// bram[9886] = 21;
// bram[9887] = 14;
// bram[9888] = 8;
// bram[9889] = 3;
// bram[9890] = 1;
// bram[9891] = 0;
// bram[9892] = 0;
// bram[9893] = 2;
// bram[9894] = 6;
// bram[9895] = 12;
// bram[9896] = 19;
// bram[9897] = 27;
// bram[9898] = 37;
// bram[9899] = 48;
// bram[9900] = 60;
// bram[9901] = 73;
// bram[9902] = 87;
// bram[9903] = 101;
// bram[9904] = 115;
// bram[9905] = 130;
// bram[9906] = 145;
// bram[9907] = 159;
// bram[9908] = 173;
// bram[9909] = 186;
// bram[9910] = 199;
// bram[9911] = 210;
// bram[9912] = 221;
// bram[9913] = 230;
// bram[9914] = 238;
// bram[9915] = 244;
// bram[9916] = 249;
// bram[9917] = 252;
// bram[9918] = 253;
// bram[9919] = 253;
// bram[9920] = 251;
// bram[9921] = 248;
// bram[9922] = 242;
// bram[9923] = 236;
// bram[9924] = 228;
// bram[9925] = 218;
// bram[9926] = 207;
// bram[9927] = 195;
// bram[9928] = 183;
// bram[9929] = 169;
// bram[9930] = 155;
// bram[9931] = 141;
// bram[9932] = 126;
// bram[9933] = 111;
// bram[9934] = 97;
// bram[9935] = 83;
// bram[9936] = 70;
// bram[9937] = 57;
// bram[9938] = 45;
// bram[9939] = 34;
// bram[9940] = 25;
// bram[9941] = 17;
// bram[9942] = 10;
// bram[9943] = 5;
// bram[9944] = 2;
// bram[9945] = 0;
// bram[9946] = 0;
// bram[9947] = 1;
// bram[9948] = 4;
// bram[9949] = 9;
// bram[9950] = 16;
// bram[9951] = 24;
// bram[9952] = 33;
// bram[9953] = 43;
// bram[9954] = 55;
// bram[9955] = 68;
// bram[9956] = 81;
// bram[9957] = 95;
// bram[9958] = 109;
// bram[9959] = 124;
// bram[9960] = 138;
// bram[9961] = 153;
// bram[9962] = 167;
// bram[9963] = 181;
// bram[9964] = 194;
// bram[9965] = 206;
// bram[9966] = 216;
// bram[9967] = 226;
// bram[9968] = 235;
// bram[9969] = 242;
// bram[9970] = 247;
// bram[9971] = 251;
// bram[9972] = 253;
// bram[9973] = 253;
// bram[9974] = 252;
// bram[9975] = 249;
// bram[9976] = 245;
// bram[9977] = 239;
// bram[9978] = 231;
// bram[9979] = 222;
// bram[9980] = 212;
// bram[9981] = 201;
// bram[9982] = 188;
// bram[9983] = 175;
// bram[9984] = 161;
// bram[9985] = 147;
// bram[9986] = 132;
// bram[9987] = 118;
// bram[9988] = 103;
// bram[9989] = 89;
// bram[9990] = 75;
// bram[9991] = 62;
// bram[9992] = 50;
// bram[9993] = 39;
// bram[9994] = 29;
// bram[9995] = 20;
// bram[9996] = 13;
// bram[9997] = 7;
// bram[9998] = 3;
// bram[9999] = 0;
// bram[10000] = 0;
// bram[10001] = 0;
// bram[10002] = 3;
// bram[10003] = 7;
// bram[10004] = 13;
// bram[10005] = 20;
// bram[10006] = 29;
// bram[10007] = 39;
// bram[10008] = 50;
// bram[10009] = 62;
// bram[10010] = 75;
// bram[10011] = 89;
// bram[10012] = 103;
// bram[10013] = 118;
// bram[10014] = 132;
// bram[10015] = 147;
// bram[10016] = 161;
// bram[10017] = 175;
// bram[10018] = 188;
// bram[10019] = 201;
// bram[10020] = 212;
// bram[10021] = 222;
// bram[10022] = 231;
// bram[10023] = 239;
// bram[10024] = 245;
// bram[10025] = 249;
// bram[10026] = 252;
// bram[10027] = 253;
// bram[10028] = 253;
// bram[10029] = 251;
// bram[10030] = 247;
// bram[10031] = 242;
// bram[10032] = 235;
// bram[10033] = 226;
// bram[10034] = 216;
// bram[10035] = 206;
// bram[10036] = 194;
// bram[10037] = 181;
// bram[10038] = 167;
// bram[10039] = 153;
// bram[10040] = 138;
// bram[10041] = 124;
// bram[10042] = 109;
// bram[10043] = 95;
// bram[10044] = 81;
// bram[10045] = 68;
// bram[10046] = 55;
// bram[10047] = 43;
// bram[10048] = 33;
// bram[10049] = 24;
// bram[10050] = 16;
// bram[10051] = 9;
// bram[10052] = 4;
// bram[10053] = 1;
// bram[10054] = 0;
// bram[10055] = 0;
// bram[10056] = 2;
// bram[10057] = 5;
// bram[10058] = 10;
// bram[10059] = 17;
// bram[10060] = 25;
// bram[10061] = 34;
// bram[10062] = 45;
// bram[10063] = 57;
// bram[10064] = 70;
// bram[10065] = 83;
// bram[10066] = 97;
// bram[10067] = 111;
// bram[10068] = 126;
// bram[10069] = 141;
// bram[10070] = 155;
// bram[10071] = 169;
// bram[10072] = 183;
// bram[10073] = 195;
// bram[10074] = 207;
// bram[10075] = 218;
// bram[10076] = 228;
// bram[10077] = 236;
// bram[10078] = 242;
// bram[10079] = 248;
// bram[10080] = 251;
// bram[10081] = 253;
// bram[10082] = 253;
// bram[10083] = 252;
// bram[10084] = 249;
// bram[10085] = 244;
// bram[10086] = 238;
// bram[10087] = 230;
// bram[10088] = 221;
// bram[10089] = 210;
// bram[10090] = 199;
// bram[10091] = 186;
// bram[10092] = 173;
// bram[10093] = 159;
// bram[10094] = 145;
// bram[10095] = 130;
// bram[10096] = 115;
// bram[10097] = 101;
// bram[10098] = 87;
// bram[10099] = 73;
// bram[10100] = 60;
// bram[10101] = 48;
// bram[10102] = 37;
// bram[10103] = 27;
// bram[10104] = 19;
// bram[10105] = 12;
// bram[10106] = 6;
// bram[10107] = 2;
// bram[10108] = 0;
// bram[10109] = 0;
// bram[10110] = 1;
// bram[10111] = 3;
// bram[10112] = 8;
// bram[10113] = 14;
// bram[10114] = 21;
// bram[10115] = 30;
// bram[10116] = 40;
// bram[10117] = 52;
// bram[10118] = 64;
// bram[10119] = 77;
// bram[10120] = 91;
// bram[10121] = 105;
// bram[10122] = 120;
// bram[10123] = 135;
// bram[10124] = 149;
// bram[10125] = 163;
// bram[10126] = 177;
// bram[10127] = 190;
// bram[10128] = 202;
// bram[10129] = 214;
// bram[10130] = 224;
// bram[10131] = 232;
// bram[10132] = 240;
// bram[10133] = 246;
// bram[10134] = 250;
// bram[10135] = 253;
// bram[10136] = 253;
// bram[10137] = 253;
// bram[10138] = 250;
// bram[10139] = 246;
// bram[10140] = 241;
// bram[10141] = 233;
// bram[10142] = 225;
// bram[10143] = 215;
// bram[10144] = 204;
// bram[10145] = 192;
// bram[10146] = 179;
// bram[10147] = 165;
// bram[10148] = 151;
// bram[10149] = 136;
// bram[10150] = 122;
// bram[10151] = 107;
// bram[10152] = 93;
// bram[10153] = 79;
// bram[10154] = 65;
// bram[10155] = 53;
// bram[10156] = 42;
// bram[10157] = 31;
// bram[10158] = 22;
// bram[10159] = 15;
// bram[10160] = 8;
// bram[10161] = 4;
// bram[10162] = 1;
// bram[10163] = 0;
// bram[10164] = 0;
// bram[10165] = 2;
// bram[10166] = 6;
// bram[10167] = 11;
// bram[10168] = 18;
// bram[10169] = 26;
// bram[10170] = 36;
// bram[10171] = 47;
// bram[10172] = 59;
// bram[10173] = 72;
// bram[10174] = 85;
// bram[10175] = 99;
// bram[10176] = 114;
// bram[10177] = 128;
// bram[10178] = 143;
// bram[10179] = 157;
// bram[10180] = 171;
// bram[10181] = 185;
// bram[10182] = 197;
// bram[10183] = 209;
// bram[10184] = 220;
// bram[10185] = 229;
// bram[10186] = 237;
// bram[10187] = 243;
// bram[10188] = 248;
// bram[10189] = 252;
// bram[10190] = 253;
// bram[10191] = 253;
// bram[10192] = 252;
// bram[10193] = 248;
// bram[10194] = 243;
// bram[10195] = 237;
// bram[10196] = 229;
// bram[10197] = 219;
// bram[10198] = 209;
// bram[10199] = 197;
// bram[10200] = 184;
// bram[10201] = 171;
// bram[10202] = 157;
// bram[10203] = 142;
// bram[10204] = 128;
// bram[10205] = 113;
// bram[10206] = 99;
// bram[10207] = 85;
// bram[10208] = 71;
// bram[10209] = 58;
// bram[10210] = 46;
// bram[10211] = 36;
// bram[10212] = 26;
// bram[10213] = 18;
// bram[10214] = 11;
// bram[10215] = 6;
// bram[10216] = 2;
// bram[10217] = 0;
// bram[10218] = 0;
// bram[10219] = 1;
// bram[10220] = 4;
// bram[10221] = 9;
// bram[10222] = 15;
// bram[10223] = 23;
// bram[10224] = 32;
// bram[10225] = 42;
// bram[10226] = 54;
// bram[10227] = 66;
// bram[10228] = 79;
// bram[10229] = 93;
// bram[10230] = 108;
// bram[10231] = 122;
// bram[10232] = 137;
// bram[10233] = 151;
// bram[10234] = 166;
// bram[10235] = 179;
// bram[10236] = 192;
// bram[10237] = 204;
// bram[10238] = 215;
// bram[10239] = 225;
// bram[10240] = 234;
// bram[10241] = 241;
// bram[10242] = 246;
// bram[10243] = 250;
// bram[10244] = 253;
// bram[10245] = 253;
// bram[10246] = 252;
// bram[10247] = 250;
// bram[10248] = 245;
// bram[10249] = 240;
// bram[10250] = 232;
// bram[10251] = 223;
// bram[10252] = 213;
// bram[10253] = 202;
// bram[10254] = 190;
// bram[10255] = 176;
// bram[10256] = 163;
// bram[10257] = 148;
// bram[10258] = 134;
// bram[10259] = 119;
// bram[10260] = 105;
// bram[10261] = 90;
// bram[10262] = 77;
// bram[10263] = 63;
// bram[10264] = 51;
// bram[10265] = 40;
// bram[10266] = 30;
// bram[10267] = 21;
// bram[10268] = 14;
// bram[10269] = 8;
// bram[10270] = 3;
// bram[10271] = 1;
// bram[10272] = 0;
// bram[10273] = 0;
// bram[10274] = 3;
// bram[10275] = 7;
// bram[10276] = 12;
// bram[10277] = 19;
// bram[10278] = 28;
// bram[10279] = 38;
// bram[10280] = 49;
// bram[10281] = 61;
// bram[10282] = 74;
// bram[10283] = 87;
// bram[10284] = 102;
// bram[10285] = 116;
// bram[10286] = 131;
// bram[10287] = 145;
// bram[10288] = 160;
// bram[10289] = 174;
// bram[10290] = 187;
// bram[10291] = 199;
// bram[10292] = 211;
// bram[10293] = 221;
// bram[10294] = 230;
// bram[10295] = 238;
// bram[10296] = 244;
// bram[10297] = 249;
// bram[10298] = 252;
// bram[10299] = 253;
// bram[10300] = 253;
// bram[10301] = 251;
// bram[10302] = 247;
// bram[10303] = 242;
// bram[10304] = 235;
// bram[10305] = 227;
// bram[10306] = 218;
// bram[10307] = 207;
// bram[10308] = 195;
// bram[10309] = 182;
// bram[10310] = 169;
// bram[10311] = 154;
// bram[10312] = 140;
// bram[10313] = 125;
// bram[10314] = 111;
// bram[10315] = 96;
// bram[10316] = 82;
// bram[10317] = 69;
// bram[10318] = 56;
// bram[10319] = 45;
// bram[10320] = 34;
// bram[10321] = 25;
// bram[10322] = 16;
// bram[10323] = 10;
// bram[10324] = 5;
// bram[10325] = 1;
// bram[10326] = 0;
// bram[10327] = 0;
// bram[10328] = 1;
// bram[10329] = 5;
// bram[10330] = 10;
// bram[10331] = 16;
// bram[10332] = 24;
// bram[10333] = 33;
// bram[10334] = 44;
// bram[10335] = 56;
// bram[10336] = 68;
// bram[10337] = 82;
// bram[10338] = 95;
// bram[10339] = 110;
// bram[10340] = 125;
// bram[10341] = 139;
// bram[10342] = 154;
// bram[10343] = 168;
// bram[10344] = 181;
// bram[10345] = 194;
// bram[10346] = 206;
// bram[10347] = 217;
// bram[10348] = 227;
// bram[10349] = 235;
// bram[10350] = 242;
// bram[10351] = 247;
// bram[10352] = 251;
// bram[10353] = 253;
// bram[10354] = 253;
// bram[10355] = 252;
// bram[10356] = 249;
// bram[10357] = 245;
// bram[10358] = 238;
// bram[10359] = 231;
// bram[10360] = 222;
// bram[10361] = 211;
// bram[10362] = 200;
// bram[10363] = 188;
// bram[10364] = 174;
// bram[10365] = 160;
// bram[10366] = 146;
// bram[10367] = 132;
// bram[10368] = 117;
// bram[10369] = 102;
// bram[10370] = 88;
// bram[10371] = 75;
// bram[10372] = 62;
// bram[10373] = 49;
// bram[10374] = 38;
// bram[10375] = 28;
// bram[10376] = 20;
// bram[10377] = 12;
// bram[10378] = 7;
// bram[10379] = 3;
// bram[10380] = 0;
// bram[10381] = 0;
// bram[10382] = 0;
// bram[10383] = 3;
// bram[10384] = 7;
// bram[10385] = 13;
// bram[10386] = 20;
// bram[10387] = 29;
// bram[10388] = 39;
// bram[10389] = 50;
// bram[10390] = 63;
// bram[10391] = 76;
// bram[10392] = 90;
// bram[10393] = 104;
// bram[10394] = 118;
// bram[10395] = 133;
// bram[10396] = 148;
// bram[10397] = 162;
// bram[10398] = 176;
// bram[10399] = 189;
// bram[10400] = 201;
// bram[10401] = 212;
// bram[10402] = 223;
// bram[10403] = 232;
// bram[10404] = 239;
// bram[10405] = 245;
// bram[10406] = 250;
// bram[10407] = 252;
// bram[10408] = 253;
// bram[10409] = 253;
// bram[10410] = 251;
// bram[10411] = 247;
// bram[10412] = 241;
// bram[10413] = 234;
// bram[10414] = 226;
// bram[10415] = 216;
// bram[10416] = 205;
// bram[10417] = 193;
// bram[10418] = 180;
// bram[10419] = 166;
// bram[10420] = 152;
// bram[10421] = 138;
// bram[10422] = 123;
// bram[10423] = 109;
// bram[10424] = 94;
// bram[10425] = 80;
// bram[10426] = 67;
// bram[10427] = 54;
// bram[10428] = 43;
// bram[10429] = 32;
// bram[10430] = 23;
// bram[10431] = 15;
// bram[10432] = 9;
// bram[10433] = 4;
// bram[10434] = 1;
// bram[10435] = 0;
// bram[10436] = 0;
// bram[10437] = 2;
// bram[10438] = 5;
// bram[10439] = 10;
// bram[10440] = 17;
// bram[10441] = 25;
// bram[10442] = 35;
// bram[10443] = 46;
// bram[10444] = 57;
// bram[10445] = 70;
// bram[10446] = 84;
// bram[10447] = 98;
// bram[10448] = 112;
// bram[10449] = 127;
// bram[10450] = 141;
// bram[10451] = 156;
// bram[10452] = 170;
// bram[10453] = 183;
// bram[10454] = 196;
// bram[10455] = 208;
// bram[10456] = 219;
// bram[10457] = 228;
// bram[10458] = 236;
// bram[10459] = 243;
// bram[10460] = 248;
// bram[10461] = 251;
// bram[10462] = 253;
// bram[10463] = 253;
// bram[10464] = 252;
// bram[10465] = 249;
// bram[10466] = 244;
// bram[10467] = 237;
// bram[10468] = 229;
// bram[10469] = 220;
// bram[10470] = 210;
// bram[10471] = 198;
// bram[10472] = 186;
// bram[10473] = 172;
// bram[10474] = 158;
// bram[10475] = 144;
// bram[10476] = 129;
// bram[10477] = 115;
// bram[10478] = 100;
// bram[10479] = 86;
// bram[10480] = 72;
// bram[10481] = 60;
// bram[10482] = 48;
// bram[10483] = 37;
// bram[10484] = 27;
// bram[10485] = 18;
// bram[10486] = 12;
// bram[10487] = 6;
// bram[10488] = 2;
// bram[10489] = 0;
// bram[10490] = 0;
// bram[10491] = 1;
// bram[10492] = 4;
// bram[10493] = 8;
// bram[10494] = 14;
// bram[10495] = 22;
// bram[10496] = 31;
// bram[10497] = 41;
// bram[10498] = 52;
// bram[10499] = 65;
// bram[10500] = 78;
// bram[10501] = 92;
// bram[10502] = 106;
// bram[10503] = 121;
// bram[10504] = 135;
// bram[10505] = 150;
// bram[10506] = 164;
// bram[10507] = 178;
// bram[10508] = 191;
// bram[10509] = 203;
// bram[10510] = 214;
// bram[10511] = 224;
// bram[10512] = 233;
// bram[10513] = 240;
// bram[10514] = 246;
// bram[10515] = 250;
// bram[10516] = 253;
// bram[10517] = 253;
// bram[10518] = 253;
// bram[10519] = 250;
// bram[10520] = 246;
// bram[10521] = 240;
// bram[10522] = 233;
// bram[10523] = 224;
// bram[10524] = 214;
// bram[10525] = 203;
// bram[10526] = 191;
// bram[10527] = 178;
// bram[10528] = 164;
// bram[10529] = 150;
// bram[10530] = 135;
// bram[10531] = 121;
// bram[10532] = 106;
// bram[10533] = 92;
// bram[10534] = 78;
// bram[10535] = 65;
// bram[10536] = 52;
// bram[10537] = 41;
// bram[10538] = 31;
// bram[10539] = 22;
// bram[10540] = 14;
// bram[10541] = 8;
// bram[10542] = 4;
// bram[10543] = 1;
// bram[10544] = 0;
// bram[10545] = 0;
// bram[10546] = 2;
// bram[10547] = 6;
// bram[10548] = 11;
// bram[10549] = 18;
// bram[10550] = 27;
// bram[10551] = 36;
// bram[10552] = 47;
// bram[10553] = 59;
// bram[10554] = 72;
// bram[10555] = 86;
// bram[10556] = 100;
// bram[10557] = 114;
// bram[10558] = 129;
// bram[10559] = 144;
// bram[10560] = 158;
// bram[10561] = 172;
// bram[10562] = 185;
// bram[10563] = 198;
// bram[10564] = 210;
// bram[10565] = 220;
// bram[10566] = 229;
// bram[10567] = 237;
// bram[10568] = 244;
// bram[10569] = 249;
// bram[10570] = 252;
// bram[10571] = 253;
// bram[10572] = 253;
// bram[10573] = 251;
// bram[10574] = 248;
// bram[10575] = 243;
// bram[10576] = 236;
// bram[10577] = 228;
// bram[10578] = 219;
// bram[10579] = 208;
// bram[10580] = 196;
// bram[10581] = 184;
// bram[10582] = 170;
// bram[10583] = 156;
// bram[10584] = 142;
// bram[10585] = 127;
// bram[10586] = 112;
// bram[10587] = 98;
// bram[10588] = 84;
// bram[10589] = 70;
// bram[10590] = 58;
// bram[10591] = 46;
// bram[10592] = 35;
// bram[10593] = 25;
// bram[10594] = 17;
// bram[10595] = 11;
// bram[10596] = 5;
// bram[10597] = 2;
// bram[10598] = 0;
// bram[10599] = 0;
// bram[10600] = 1;
// bram[10601] = 4;
// bram[10602] = 9;
// bram[10603] = 15;
// bram[10604] = 23;
// bram[10605] = 32;
// bram[10606] = 43;
// bram[10607] = 54;
// bram[10608] = 67;
// bram[10609] = 80;
// bram[10610] = 94;
// bram[10611] = 108;
// bram[10612] = 123;
// bram[10613] = 138;
// bram[10614] = 152;
// bram[10615] = 166;
// bram[10616] = 180;
// bram[10617] = 193;
// bram[10618] = 205;
// bram[10619] = 216;
// bram[10620] = 226;
// bram[10621] = 234;
// bram[10622] = 241;
// bram[10623] = 247;
// bram[10624] = 251;
// bram[10625] = 253;
// bram[10626] = 253;
// bram[10627] = 252;
// bram[10628] = 250;
// bram[10629] = 245;
// bram[10630] = 239;
// bram[10631] = 232;
// bram[10632] = 223;
// bram[10633] = 213;
// bram[10634] = 201;
// bram[10635] = 189;
// bram[10636] = 176;
// bram[10637] = 162;
// bram[10638] = 148;
// bram[10639] = 133;
// bram[10640] = 119;
// bram[10641] = 104;
// bram[10642] = 90;
// bram[10643] = 76;
// bram[10644] = 63;
// bram[10645] = 51;
// bram[10646] = 39;
// bram[10647] = 29;
// bram[10648] = 21;
// bram[10649] = 13;
// bram[10650] = 7;
// bram[10651] = 3;
// bram[10652] = 0;
// bram[10653] = 0;
// bram[10654] = 0;
// bram[10655] = 3;
// bram[10656] = 7;
// bram[10657] = 12;
// bram[10658] = 20;
// bram[10659] = 28;
// bram[10660] = 38;
// bram[10661] = 49;
// bram[10662] = 61;
// bram[10663] = 74;
// bram[10664] = 88;
// bram[10665] = 102;
// bram[10666] = 117;
// bram[10667] = 131;
// bram[10668] = 146;
// bram[10669] = 160;
// bram[10670] = 174;
// bram[10671] = 187;
// bram[10672] = 200;
// bram[10673] = 211;
// bram[10674] = 222;
// bram[10675] = 231;
// bram[10676] = 238;
// bram[10677] = 245;
// bram[10678] = 249;
// bram[10679] = 252;
// bram[10680] = 253;
// bram[10681] = 253;
// bram[10682] = 251;
// bram[10683] = 247;
// bram[10684] = 242;
// bram[10685] = 235;
// bram[10686] = 227;
// bram[10687] = 217;
// bram[10688] = 206;
// bram[10689] = 194;
// bram[10690] = 181;
// bram[10691] = 168;
// bram[10692] = 154;
// bram[10693] = 139;
// bram[10694] = 125;
// bram[10695] = 110;
// bram[10696] = 96;
// bram[10697] = 82;
// bram[10698] = 68;
// bram[10699] = 56;
// bram[10700] = 44;
// bram[10701] = 33;
// bram[10702] = 24;
// bram[10703] = 16;
// bram[10704] = 10;
// bram[10705] = 5;
// bram[10706] = 1;
// bram[10707] = 0;
// bram[10708] = 0;
// bram[10709] = 1;
// bram[10710] = 5;
// bram[10711] = 10;
// bram[10712] = 16;
// bram[10713] = 24;
// bram[10714] = 34;
// bram[10715] = 44;
// bram[10716] = 56;
// bram[10717] = 69;
// bram[10718] = 82;
// bram[10719] = 96;
// bram[10720] = 111;
// bram[10721] = 125;
// bram[10722] = 140;
// bram[10723] = 154;
// bram[10724] = 168;
// bram[10725] = 182;
// bram[10726] = 195;
// bram[10727] = 207;
// bram[10728] = 217;
// bram[10729] = 227;
// bram[10730] = 235;
// bram[10731] = 242;
// bram[10732] = 247;
// bram[10733] = 251;
// bram[10734] = 253;
// bram[10735] = 253;
// bram[10736] = 252;
// bram[10737] = 249;
// bram[10738] = 244;
// bram[10739] = 238;
// bram[10740] = 230;
// bram[10741] = 221;
// bram[10742] = 211;
// bram[10743] = 199;
// bram[10744] = 187;
// bram[10745] = 174;
// bram[10746] = 160;
// bram[10747] = 145;
// bram[10748] = 131;
// bram[10749] = 116;
// bram[10750] = 102;
// bram[10751] = 88;
// bram[10752] = 74;
// bram[10753] = 61;
// bram[10754] = 49;
// bram[10755] = 38;
// bram[10756] = 28;
// bram[10757] = 19;
// bram[10758] = 12;
// bram[10759] = 7;
// bram[10760] = 3;
// bram[10761] = 0;
// bram[10762] = 0;
// bram[10763] = 1;
// bram[10764] = 3;
// bram[10765] = 8;
// bram[10766] = 13;
// bram[10767] = 21;
// bram[10768] = 30;
// bram[10769] = 40;
// bram[10770] = 51;
// bram[10771] = 63;
// bram[10772] = 76;
// bram[10773] = 90;
// bram[10774] = 104;
// bram[10775] = 119;
// bram[10776] = 134;
// bram[10777] = 148;
// bram[10778] = 163;
// bram[10779] = 176;
// bram[10780] = 189;
// bram[10781] = 202;
// bram[10782] = 213;
// bram[10783] = 223;
// bram[10784] = 232;
// bram[10785] = 239;
// bram[10786] = 245;
// bram[10787] = 250;
// bram[10788] = 252;
// bram[10789] = 253;
// bram[10790] = 253;
// bram[10791] = 251;
// bram[10792] = 247;
// bram[10793] = 241;
// bram[10794] = 234;
// bram[10795] = 225;
// bram[10796] = 215;
// bram[10797] = 204;
// bram[10798] = 192;
// bram[10799] = 179;
// bram[10800] = 166;
// bram[10801] = 152;
// bram[10802] = 137;
// bram[10803] = 122;
// bram[10804] = 108;
// bram[10805] = 93;
// bram[10806] = 80;
// bram[10807] = 66;
// bram[10808] = 54;
// bram[10809] = 42;
// bram[10810] = 32;
// bram[10811] = 23;
// bram[10812] = 15;
// bram[10813] = 9;
// bram[10814] = 4;
// bram[10815] = 1;
// bram[10816] = 0;
// bram[10817] = 0;
// bram[10818] = 2;
// bram[10819] = 6;
// bram[10820] = 11;
// bram[10821] = 18;
// bram[10822] = 26;
// bram[10823] = 35;
// bram[10824] = 46;
// bram[10825] = 58;
// bram[10826] = 71;
// bram[10827] = 84;
// bram[10828] = 98;
// bram[10829] = 113;
// bram[10830] = 127;
// bram[10831] = 142;
// bram[10832] = 157;
// bram[10833] = 171;
// bram[10834] = 184;
// bram[10835] = 197;
// bram[10836] = 208;
// bram[10837] = 219;
// bram[10838] = 228;
// bram[10839] = 236;
// bram[10840] = 243;
// bram[10841] = 248;
// bram[10842] = 252;
// bram[10843] = 253;
// bram[10844] = 253;
// bram[10845] = 252;
// bram[10846] = 248;
// bram[10847] = 243;
// bram[10848] = 237;
// bram[10849] = 229;
// bram[10850] = 220;
// bram[10851] = 209;
// bram[10852] = 198;
// bram[10853] = 185;
// bram[10854] = 172;
// bram[10855] = 158;
// bram[10856] = 143;
// bram[10857] = 129;
// bram[10858] = 114;
// bram[10859] = 99;
// bram[10860] = 85;
// bram[10861] = 72;
// bram[10862] = 59;
// bram[10863] = 47;
// bram[10864] = 36;
// bram[10865] = 26;
// bram[10866] = 18;
// bram[10867] = 11;
// bram[10868] = 6;
// bram[10869] = 2;
// bram[10870] = 0;
// bram[10871] = 0;
// bram[10872] = 1;
// bram[10873] = 4;
// bram[10874] = 8;
// bram[10875] = 14;
// bram[10876] = 22;
// bram[10877] = 31;
// bram[10878] = 41;
// bram[10879] = 53;
// bram[10880] = 65;
// bram[10881] = 79;
// bram[10882] = 92;
// bram[10883] = 107;
// bram[10884] = 121;
// bram[10885] = 136;
// bram[10886] = 150;
// bram[10887] = 165;
// bram[10888] = 178;
// bram[10889] = 191;
// bram[10890] = 204;
// bram[10891] = 215;
// bram[10892] = 225;
// bram[10893] = 233;
// bram[10894] = 240;
// bram[10895] = 246;
// bram[10896] = 250;
// bram[10897] = 253;
// bram[10898] = 253;
// bram[10899] = 253;
// bram[10900] = 250;
// bram[10901] = 246;
// bram[10902] = 240;
// bram[10903] = 233;
// bram[10904] = 224;
// bram[10905] = 214;
// bram[10906] = 203;
// bram[10907] = 190;
// bram[10908] = 177;
// bram[10909] = 164;
// bram[10910] = 149;
// bram[10911] = 135;
// bram[10912] = 120;
// bram[10913] = 106;
// bram[10914] = 91;
// bram[10915] = 77;
// bram[10916] = 64;
// bram[10917] = 52;
// bram[10918] = 41;
// bram[10919] = 30;
// bram[10920] = 21;
// bram[10921] = 14;
// bram[10922] = 8;
// bram[10923] = 3;
// bram[10924] = 1;
// bram[10925] = 0;
// bram[10926] = 0;
// bram[10927] = 2;
// bram[10928] = 6;
// bram[10929] = 12;
// bram[10930] = 19;
// bram[10931] = 27;
// bram[10932] = 37;
// bram[10933] = 48;
// bram[10934] = 60;
// bram[10935] = 73;
// bram[10936] = 86;
// bram[10937] = 101;
// bram[10938] = 115;
// bram[10939] = 130;
// bram[10940] = 144;
// bram[10941] = 159;
// bram[10942] = 173;
// bram[10943] = 186;
// bram[10944] = 199;
// bram[10945] = 210;
// bram[10946] = 221;
// bram[10947] = 230;
// bram[10948] = 238;
// bram[10949] = 244;
// bram[10950] = 249;
// bram[10951] = 252;
// bram[10952] = 253;
// bram[10953] = 253;
// bram[10954] = 251;
// bram[10955] = 248;
// bram[10956] = 243;
// bram[10957] = 236;
// bram[10958] = 228;
// bram[10959] = 218;
// bram[10960] = 207;
// bram[10961] = 196;
// bram[10962] = 183;
// bram[10963] = 169;
// bram[10964] = 155;
// bram[10965] = 141;
// bram[10966] = 126;
// bram[10967] = 112;
// bram[10968] = 97;
// bram[10969] = 83;
// bram[10970] = 70;
// bram[10971] = 57;
// bram[10972] = 45;
// bram[10973] = 35;
// bram[10974] = 25;
// bram[10975] = 17;
// bram[10976] = 10;
// bram[10977] = 5;
// bram[10978] = 2;
// bram[10979] = 0;
// bram[10980] = 0;
// bram[10981] = 1;
// bram[10982] = 4;
// bram[10983] = 9;
// bram[10984] = 16;
// bram[10985] = 23;
// bram[10986] = 33;
// bram[10987] = 43;
// bram[10988] = 55;
// bram[10989] = 67;
// bram[10990] = 81;
// bram[10991] = 95;
// bram[10992] = 109;
// bram[10993] = 124;
// bram[10994] = 138;
// bram[10995] = 153;
// bram[10996] = 167;
// bram[10997] = 180;
// bram[10998] = 193;
// bram[10999] = 205;
// bram[11000] = 216;
// bram[11001] = 226;
// bram[11002] = 234;
// bram[11003] = 241;
// bram[11004] = 247;
// bram[11005] = 251;
// bram[11006] = 253;
// bram[11007] = 253;
// bram[11008] = 252;
// bram[11009] = 249;
// bram[11010] = 245;
// bram[11011] = 239;
// bram[11012] = 231;
// bram[11013] = 222;
// bram[11014] = 212;
// bram[11015] = 201;
// bram[11016] = 188;
// bram[11017] = 175;
// bram[11018] = 161;
// bram[11019] = 147;
// bram[11020] = 132;
// bram[11021] = 118;
// bram[11022] = 103;
// bram[11023] = 89;
// bram[11024] = 75;
// bram[11025] = 62;
// bram[11026] = 50;
// bram[11027] = 39;
// bram[11028] = 29;
// bram[11029] = 20;
// bram[11030] = 13;
// bram[11031] = 7;
// bram[11032] = 3;
// bram[11033] = 0;
// bram[11034] = 0;
// bram[11035] = 0;
// bram[11036] = 3;
// bram[11037] = 7;
// bram[11038] = 13;
// bram[11039] = 20;
// bram[11040] = 29;
// bram[11041] = 39;
// bram[11042] = 50;
// bram[11043] = 62;
// bram[11044] = 75;
// bram[11045] = 89;
// bram[11046] = 103;
// bram[11047] = 117;
// bram[11048] = 132;
// bram[11049] = 147;
// bram[11050] = 161;
// bram[11051] = 175;
// bram[11052] = 188;
// bram[11053] = 200;
// bram[11054] = 212;
// bram[11055] = 222;
// bram[11056] = 231;
// bram[11057] = 239;
// bram[11058] = 245;
// bram[11059] = 249;
// bram[11060] = 252;
// bram[11061] = 253;
// bram[11062] = 253;
// bram[11063] = 251;
// bram[11064] = 247;
// bram[11065] = 242;
// bram[11066] = 235;
// bram[11067] = 226;
// bram[11068] = 217;
// bram[11069] = 206;
// bram[11070] = 194;
// bram[11071] = 181;
// bram[11072] = 167;
// bram[11073] = 153;
// bram[11074] = 139;
// bram[11075] = 124;
// bram[11076] = 109;
// bram[11077] = 95;
// bram[11078] = 81;
// bram[11079] = 68;
// bram[11080] = 55;
// bram[11081] = 43;
// bram[11082] = 33;
// bram[11083] = 24;
// bram[11084] = 16;
// bram[11085] = 9;
// bram[11086] = 4;
// bram[11087] = 1;
// bram[11088] = 0;
// bram[11089] = 0;
// bram[11090] = 2;
// bram[11091] = 5;
// bram[11092] = 10;
// bram[11093] = 17;
// bram[11094] = 25;
// bram[11095] = 34;
// bram[11096] = 45;
// bram[11097] = 57;
// bram[11098] = 69;
// bram[11099] = 83;
// bram[11100] = 97;
// bram[11101] = 111;
// bram[11102] = 126;
// bram[11103] = 141;
// bram[11104] = 155;
// bram[11105] = 169;
// bram[11106] = 183;
// bram[11107] = 195;
// bram[11108] = 207;
// bram[11109] = 218;
// bram[11110] = 227;
// bram[11111] = 236;
// bram[11112] = 242;
// bram[11113] = 248;
// bram[11114] = 251;
// bram[11115] = 253;
// bram[11116] = 253;
// bram[11117] = 252;
// bram[11118] = 249;
// bram[11119] = 244;
// bram[11120] = 238;
// bram[11121] = 230;
// bram[11122] = 221;
// bram[11123] = 210;
// bram[11124] = 199;
// bram[11125] = 186;
// bram[11126] = 173;
// bram[11127] = 159;
// bram[11128] = 145;
// bram[11129] = 130;
// bram[11130] = 116;
// bram[11131] = 101;
// bram[11132] = 87;
// bram[11133] = 73;
// bram[11134] = 60;
// bram[11135] = 48;
// bram[11136] = 37;
// bram[11137] = 27;
// bram[11138] = 19;
// bram[11139] = 12;
// bram[11140] = 6;
// bram[11141] = 2;
// bram[11142] = 0;
// bram[11143] = 0;
// bram[11144] = 1;
// bram[11145] = 3;
// bram[11146] = 8;
// bram[11147] = 14;
// bram[11148] = 21;
// bram[11149] = 30;
// bram[11150] = 40;
// bram[11151] = 52;
// bram[11152] = 64;
// bram[11153] = 77;
// bram[11154] = 91;
// bram[11155] = 105;
// bram[11156] = 120;
// bram[11157] = 134;
// bram[11158] = 149;
// bram[11159] = 163;
// bram[11160] = 177;
// bram[11161] = 190;
// bram[11162] = 202;
// bram[11163] = 214;
// bram[11164] = 224;
// bram[11165] = 232;
// bram[11166] = 240;
// bram[11167] = 246;
// bram[11168] = 250;
// bram[11169] = 253;
// bram[11170] = 253;
// bram[11171] = 253;
// bram[11172] = 250;
// bram[11173] = 246;
// bram[11174] = 241;
// bram[11175] = 233;
// bram[11176] = 225;
// bram[11177] = 215;
// bram[11178] = 204;
// bram[11179] = 192;
// bram[11180] = 179;
// bram[11181] = 165;
// bram[11182] = 151;
// bram[11183] = 136;
// bram[11184] = 122;
// bram[11185] = 107;
// bram[11186] = 93;
// bram[11187] = 79;
// bram[11188] = 66;
// bram[11189] = 53;
// bram[11190] = 42;
// bram[11191] = 31;
// bram[11192] = 22;
// bram[11193] = 15;
// bram[11194] = 8;
// bram[11195] = 4;
// bram[11196] = 1;
// bram[11197] = 0;
// bram[11198] = 0;
// bram[11199] = 2;
// bram[11200] = 6;
// bram[11201] = 11;
// bram[11202] = 18;
// bram[11203] = 26;
// bram[11204] = 36;
// bram[11205] = 47;
// bram[11206] = 59;
// bram[11207] = 71;
// bram[11208] = 85;
// bram[11209] = 99;
// bram[11210] = 114;
// bram[11211] = 128;
// bram[11212] = 143;
// bram[11213] = 157;
// bram[11214] = 171;
// bram[11215] = 185;
// bram[11216] = 197;
// bram[11217] = 209;
// bram[11218] = 219;
// bram[11219] = 229;
// bram[11220] = 237;
// bram[11221] = 243;
// bram[11222] = 248;
// bram[11223] = 252;
// bram[11224] = 253;
// bram[11225] = 253;
// bram[11226] = 252;
// bram[11227] = 248;
// bram[11228] = 243;
// bram[11229] = 237;
// bram[11230] = 229;
// bram[11231] = 219;
// bram[11232] = 209;
// bram[11233] = 197;
// bram[11234] = 184;
// bram[11235] = 171;
// bram[11236] = 157;
// bram[11237] = 143;
// bram[11238] = 128;
// bram[11239] = 113;
// bram[11240] = 99;
// bram[11241] = 85;
// bram[11242] = 71;
// bram[11243] = 58;
// bram[11244] = 46;
// bram[11245] = 36;
// bram[11246] = 26;
// bram[11247] = 18;
// bram[11248] = 11;
// bram[11249] = 6;
// bram[11250] = 2;
// bram[11251] = 0;
// bram[11252] = 0;
// bram[11253] = 1;
// bram[11254] = 4;
// bram[11255] = 9;
// bram[11256] = 15;
// bram[11257] = 23;
// bram[11258] = 32;
// bram[11259] = 42;
// bram[11260] = 53;
// bram[11261] = 66;
// bram[11262] = 79;
// bram[11263] = 93;
// bram[11264] = 107;
// bram[11265] = 122;
// bram[11266] = 137;
// bram[11267] = 151;
// bram[11268] = 165;
// bram[11269] = 179;
// bram[11270] = 192;
// bram[11271] = 204;
// bram[11272] = 215;
// bram[11273] = 225;
// bram[11274] = 234;
// bram[11275] = 241;
// bram[11276] = 246;
// bram[11277] = 250;
// bram[11278] = 253;
// bram[11279] = 253;
// bram[11280] = 252;
// bram[11281] = 250;
// bram[11282] = 246;
// bram[11283] = 240;
// bram[11284] = 232;
// bram[11285] = 223;
// bram[11286] = 213;
// bram[11287] = 202;
// bram[11288] = 190;
// bram[11289] = 177;
// bram[11290] = 163;
// bram[11291] = 149;
// bram[11292] = 134;
// bram[11293] = 119;
// bram[11294] = 105;
// bram[11295] = 91;
// bram[11296] = 77;
// bram[11297] = 64;
// bram[11298] = 51;
// bram[11299] = 40;
// bram[11300] = 30;
// bram[11301] = 21;
// bram[11302] = 14;
// bram[11303] = 8;
// bram[11304] = 3;
// bram[11305] = 1;
// bram[11306] = 0;
// bram[11307] = 0;
// bram[11308] = 2;
// bram[11309] = 6;
// bram[11310] = 12;
// bram[11311] = 19;
// bram[11312] = 28;
// bram[11313] = 37;
// bram[11314] = 49;
// bram[11315] = 61;
// bram[11316] = 74;
// bram[11317] = 87;
// bram[11318] = 101;
// bram[11319] = 116;
// bram[11320] = 130;
// bram[11321] = 145;
// bram[11322] = 159;
// bram[11323] = 173;
// bram[11324] = 187;
// bram[11325] = 199;
// bram[11326] = 211;
// bram[11327] = 221;
// bram[11328] = 230;
// bram[11329] = 238;
// bram[11330] = 244;
// bram[11331] = 249;
// bram[11332] = 252;
// bram[11333] = 253;
// bram[11334] = 253;
// bram[11335] = 251;
// bram[11336] = 248;
// bram[11337] = 242;
// bram[11338] = 236;
// bram[11339] = 227;
// bram[11340] = 218;
// bram[11341] = 207;
// bram[11342] = 195;
// bram[11343] = 182;
// bram[11344] = 169;
// bram[11345] = 155;
// bram[11346] = 140;
// bram[11347] = 126;
// bram[11348] = 111;
// bram[11349] = 97;
// bram[11350] = 83;
// bram[11351] = 69;
// bram[11352] = 56;
// bram[11353] = 45;
// bram[11354] = 34;
// bram[11355] = 25;
// bram[11356] = 17;
// bram[11357] = 10;
// bram[11358] = 5;
// bram[11359] = 2;
// bram[11360] = 0;
// bram[11361] = 0;
// bram[11362] = 1;
// bram[11363] = 5;
// bram[11364] = 9;
// bram[11365] = 16;
// bram[11366] = 24;
// bram[11367] = 33;
// bram[11368] = 44;
// bram[11369] = 55;
// bram[11370] = 68;
// bram[11371] = 81;
// bram[11372] = 95;
// bram[11373] = 110;
// bram[11374] = 124;
// bram[11375] = 139;
// bram[11376] = 153;
// bram[11377] = 168;
// bram[11378] = 181;
// bram[11379] = 194;
// bram[11380] = 206;
// bram[11381] = 217;
// bram[11382] = 226;
// bram[11383] = 235;
// bram[11384] = 242;
// bram[11385] = 247;
// bram[11386] = 251;
// bram[11387] = 253;
// bram[11388] = 253;
// bram[11389] = 252;
// bram[11390] = 249;
// bram[11391] = 245;
// bram[11392] = 239;
// bram[11393] = 231;
// bram[11394] = 222;
// bram[11395] = 212;
// bram[11396] = 200;
// bram[11397] = 188;
// bram[11398] = 175;
// bram[11399] = 161;
// bram[11400] = 146;
// bram[11401] = 132;
// bram[11402] = 117;
// bram[11403] = 103;
// bram[11404] = 88;
// bram[11405] = 75;
// bram[11406] = 62;
// bram[11407] = 50;
// bram[11408] = 38;
// bram[11409] = 28;
// bram[11410] = 20;
// bram[11411] = 13;
// bram[11412] = 7;
// bram[11413] = 3;
// bram[11414] = 0;
// bram[11415] = 0;
// bram[11416] = 0;
// bram[11417] = 3;
// bram[11418] = 7;
// bram[11419] = 13;
// bram[11420] = 20;
// bram[11421] = 29;
// bram[11422] = 39;
// bram[11423] = 50;
// bram[11424] = 63;
// bram[11425] = 76;
// bram[11426] = 89;
// bram[11427] = 104;
// bram[11428] = 118;
// bram[11429] = 133;
// bram[11430] = 147;
// bram[11431] = 162;
// bram[11432] = 175;
// bram[11433] = 189;
// bram[11434] = 201;
// bram[11435] = 212;
// bram[11436] = 223;
// bram[11437] = 231;
// bram[11438] = 239;
// bram[11439] = 245;
// bram[11440] = 250;
// bram[11441] = 252;
// bram[11442] = 253;
// bram[11443] = 253;
// bram[11444] = 251;
// bram[11445] = 247;
// bram[11446] = 241;
// bram[11447] = 234;
// bram[11448] = 226;
// bram[11449] = 216;
// bram[11450] = 205;
// bram[11451] = 193;
// bram[11452] = 180;
// bram[11453] = 167;
// bram[11454] = 152;
// bram[11455] = 138;
// bram[11456] = 123;
// bram[11457] = 109;
// bram[11458] = 94;
// bram[11459] = 80;
// bram[11460] = 67;
// bram[11461] = 55;
// bram[11462] = 43;
// bram[11463] = 32;
// bram[11464] = 23;
// bram[11465] = 15;
// bram[11466] = 9;
// bram[11467] = 4;
// bram[11468] = 1;
// bram[11469] = 0;
// bram[11470] = 0;
// bram[11471] = 2;
// bram[11472] = 5;
// bram[11473] = 10;
// bram[11474] = 17;
// bram[11475] = 25;
// bram[11476] = 35;
// bram[11477] = 45;
// bram[11478] = 57;
// bram[11479] = 70;
// bram[11480] = 83;
// bram[11481] = 98;
// bram[11482] = 112;
// bram[11483] = 127;
// bram[11484] = 141;
// bram[11485] = 156;
// bram[11486] = 170;
// bram[11487] = 183;
// bram[11488] = 196;
// bram[11489] = 208;
// bram[11490] = 218;
// bram[11491] = 228;
// bram[11492] = 236;
// bram[11493] = 243;
// bram[11494] = 248;
// bram[11495] = 251;
// bram[11496] = 253;
// bram[11497] = 253;
// bram[11498] = 252;
// bram[11499] = 249;
// bram[11500] = 244;
// bram[11501] = 237;
// bram[11502] = 230;
// bram[11503] = 220;
// bram[11504] = 210;
// bram[11505] = 198;
// bram[11506] = 186;
// bram[11507] = 172;
// bram[11508] = 158;
// bram[11509] = 144;
// bram[11510] = 129;
// bram[11511] = 115;
// bram[11512] = 100;
// bram[11513] = 86;
// bram[11514] = 73;
// bram[11515] = 60;
// bram[11516] = 48;
// bram[11517] = 37;
// bram[11518] = 27;
// bram[11519] = 19;
// bram[11520] = 12;
// bram[11521] = 6;
// bram[11522] = 2;
// bram[11523] = 0;
// bram[11524] = 0;
// bram[11525] = 1;
// bram[11526] = 4;
// bram[11527] = 8;
// bram[11528] = 14;
// bram[11529] = 22;
// bram[11530] = 31;
// bram[11531] = 41;
// bram[11532] = 52;
// bram[11533] = 65;
// bram[11534] = 78;
// bram[11535] = 92;
// bram[11536] = 106;
// bram[11537] = 120;
// bram[11538] = 135;
// bram[11539] = 150;
// bram[11540] = 164;
// bram[11541] = 178;
// bram[11542] = 191;
// bram[11543] = 203;
// bram[11544] = 214;
// bram[11545] = 224;
// bram[11546] = 233;
// bram[11547] = 240;
// bram[11548] = 246;
// bram[11549] = 250;
// bram[11550] = 253;
// bram[11551] = 253;
// bram[11552] = 253;
// bram[11553] = 250;
// bram[11554] = 246;
// bram[11555] = 240;
// bram[11556] = 233;
// bram[11557] = 224;
// bram[11558] = 214;
// bram[11559] = 203;
// bram[11560] = 191;
// bram[11561] = 178;
// bram[11562] = 164;
// bram[11563] = 150;
// bram[11564] = 136;
// bram[11565] = 121;
// bram[11566] = 106;
// bram[11567] = 92;
// bram[11568] = 78;
// bram[11569] = 65;
// bram[11570] = 53;
// bram[11571] = 41;
// bram[11572] = 31;
// bram[11573] = 22;
// bram[11574] = 14;
// bram[11575] = 8;
// bram[11576] = 4;
// bram[11577] = 1;
// bram[11578] = 0;
// bram[11579] = 0;
// bram[11580] = 2;
// bram[11581] = 6;
// bram[11582] = 11;
// bram[11583] = 18;
// bram[11584] = 27;
// bram[11585] = 36;
// bram[11586] = 47;
// bram[11587] = 59;
// bram[11588] = 72;
// bram[11589] = 86;
// bram[11590] = 100;
// bram[11591] = 114;
// bram[11592] = 129;
// bram[11593] = 144;
// bram[11594] = 158;
// bram[11595] = 172;
// bram[11596] = 185;
// bram[11597] = 198;
// bram[11598] = 209;
// bram[11599] = 220;
// bram[11600] = 229;
// bram[11601] = 237;
// bram[11602] = 244;
// bram[11603] = 248;
// bram[11604] = 252;
// bram[11605] = 253;
// bram[11606] = 253;
// bram[11607] = 251;
// bram[11608] = 248;
// bram[11609] = 243;
// bram[11610] = 236;
// bram[11611] = 228;
// bram[11612] = 219;
// bram[11613] = 208;
// bram[11614] = 196;
// bram[11615] = 184;
// bram[11616] = 170;
// bram[11617] = 156;
// bram[11618] = 142;
// bram[11619] = 127;
// bram[11620] = 113;
// bram[11621] = 98;
// bram[11622] = 84;
// bram[11623] = 71;
// bram[11624] = 58;
// bram[11625] = 46;
// bram[11626] = 35;
// bram[11627] = 26;
// bram[11628] = 17;
// bram[11629] = 11;
// bram[11630] = 5;
// bram[11631] = 2;
// bram[11632] = 0;
// bram[11633] = 0;
// bram[11634] = 1;
// bram[11635] = 4;
// bram[11636] = 9;
// bram[11637] = 15;
// bram[11638] = 23;
// bram[11639] = 32;
// bram[11640] = 43;
// bram[11641] = 54;
// bram[11642] = 67;
// bram[11643] = 80;
// bram[11644] = 94;
// bram[11645] = 108;
// bram[11646] = 123;
// bram[11647] = 137;
// bram[11648] = 152;
// bram[11649] = 166;
// bram[11650] = 180;
// bram[11651] = 193;
// bram[11652] = 205;
// bram[11653] = 216;
// bram[11654] = 225;
// bram[11655] = 234;
// bram[11656] = 241;
// bram[11657] = 247;
// bram[11658] = 251;
// bram[11659] = 253;
// bram[11660] = 253;
// bram[11661] = 252;
// bram[11662] = 250;
// bram[11663] = 245;
// bram[11664] = 239;
// bram[11665] = 232;
// bram[11666] = 223;
// bram[11667] = 213;
// bram[11668] = 201;
// bram[11669] = 189;
// bram[11670] = 176;
// bram[11671] = 162;
// bram[11672] = 148;
// bram[11673] = 133;
// bram[11674] = 119;
// bram[11675] = 104;
// bram[11676] = 90;
// bram[11677] = 76;
// bram[11678] = 63;
// bram[11679] = 51;
// bram[11680] = 40;
// bram[11681] = 29;
// bram[11682] = 21;
// bram[11683] = 13;
// bram[11684] = 7;
// bram[11685] = 3;
// bram[11686] = 0;
// bram[11687] = 0;
// bram[11688] = 0;
// bram[11689] = 3;
// bram[11690] = 7;
// bram[11691] = 12;
// bram[11692] = 19;
// bram[11693] = 28;
// bram[11694] = 38;
// bram[11695] = 49;
// bram[11696] = 61;
// bram[11697] = 74;
// bram[11698] = 88;
// bram[11699] = 102;
// bram[11700] = 117;
// bram[11701] = 131;
// bram[11702] = 146;
// bram[11703] = 160;
// bram[11704] = 174;
// bram[11705] = 187;
// bram[11706] = 200;
// bram[11707] = 211;
// bram[11708] = 221;
// bram[11709] = 231;
// bram[11710] = 238;
// bram[11711] = 244;
// bram[11712] = 249;
// bram[11713] = 252;
// bram[11714] = 253;
// bram[11715] = 253;
// bram[11716] = 251;
// bram[11717] = 247;
// bram[11718] = 242;
// bram[11719] = 235;
// bram[11720] = 227;
// bram[11721] = 217;
// bram[11722] = 206;
// bram[11723] = 194;
// bram[11724] = 182;
// bram[11725] = 168;
// bram[11726] = 154;
// bram[11727] = 140;
// bram[11728] = 125;
// bram[11729] = 110;
// bram[11730] = 96;
// bram[11731] = 82;
// bram[11732] = 68;
// bram[11733] = 56;
// bram[11734] = 44;
// bram[11735] = 34;
// bram[11736] = 24;
// bram[11737] = 16;
// bram[11738] = 10;
// bram[11739] = 5;
// bram[11740] = 1;
// bram[11741] = 0;
// bram[11742] = 0;
// bram[11743] = 1;
// bram[11744] = 5;
// bram[11745] = 10;
// bram[11746] = 16;
// bram[11747] = 24;
// bram[11748] = 34;
// bram[11749] = 44;
// bram[11750] = 56;
// bram[11751] = 69;
// bram[11752] = 82;
// bram[11753] = 96;
// bram[11754] = 110;
// bram[11755] = 125;
// bram[11756] = 140;
// bram[11757] = 154;
// bram[11758] = 168;
// bram[11759] = 182;
// bram[11760] = 195;
// bram[11761] = 206;
// bram[11762] = 217;
// bram[11763] = 227;
// bram[11764] = 235;
// bram[11765] = 242;
// bram[11766] = 247;
// bram[11767] = 251;
// bram[11768] = 253;
// bram[11769] = 253;
// bram[11770] = 252;
// bram[11771] = 249;
// bram[11772] = 244;
// bram[11773] = 238;
// bram[11774] = 231;
// bram[11775] = 221;
// bram[11776] = 211;
// bram[11777] = 200;
// bram[11778] = 187;
// bram[11779] = 174;
// bram[11780] = 160;
// bram[11781] = 146;
// bram[11782] = 131;
// bram[11783] = 116;
// bram[11784] = 102;
// bram[11785] = 88;
// bram[11786] = 74;
// bram[11787] = 61;
// bram[11788] = 49;
// bram[11789] = 38;
// bram[11790] = 28;
// bram[11791] = 19;
// bram[11792] = 12;
// bram[11793] = 7;
// bram[11794] = 3;
// bram[11795] = 0;
// bram[11796] = 0;
// bram[11797] = 0;
// bram[11798] = 3;
// bram[11799] = 7;
// bram[11800] = 13;
// bram[11801] = 21;
// bram[11802] = 30;
// bram[11803] = 40;
// bram[11804] = 51;
// bram[11805] = 63;
// bram[11806] = 76;
// bram[11807] = 90;
// bram[11808] = 104;
// bram[11809] = 119;
// bram[11810] = 133;
// bram[11811] = 148;
// bram[11812] = 162;
// bram[11813] = 176;
// bram[11814] = 189;
// bram[11815] = 202;
// bram[11816] = 213;
// bram[11817] = 223;
// bram[11818] = 232;
// bram[11819] = 239;
// bram[11820] = 245;
// bram[11821] = 250;
// bram[11822] = 252;
// bram[11823] = 253;
// bram[11824] = 253;
// bram[11825] = 251;
// bram[11826] = 247;
// bram[11827] = 241;
// bram[11828] = 234;
// bram[11829] = 225;
// bram[11830] = 216;
// bram[11831] = 205;
// bram[11832] = 193;
// bram[11833] = 180;
// bram[11834] = 166;
// bram[11835] = 152;
// bram[11836] = 137;
// bram[11837] = 123;
// bram[11838] = 108;
// bram[11839] = 94;
// bram[11840] = 80;
// bram[11841] = 66;
// bram[11842] = 54;
// bram[11843] = 42;
// bram[11844] = 32;
// bram[11845] = 23;
// bram[11846] = 15;
// bram[11847] = 9;
// bram[11848] = 4;
// bram[11849] = 1;
// bram[11850] = 0;
// bram[11851] = 0;
// bram[11852] = 2;
// bram[11853] = 5;
// bram[11854] = 11;
// bram[11855] = 17;
// bram[11856] = 26;
// bram[11857] = 35;
// bram[11858] = 46;
// bram[11859] = 58;
// bram[11860] = 71;
// bram[11861] = 84;
// bram[11862] = 98;
// bram[11863] = 113;
// bram[11864] = 127;
// bram[11865] = 142;
// bram[11866] = 156;
// bram[11867] = 170;
// bram[11868] = 184;
// bram[11869] = 196;
// bram[11870] = 208;
// bram[11871] = 219;
// bram[11872] = 228;
// bram[11873] = 236;
// bram[11874] = 243;
// bram[11875] = 248;
// bram[11876] = 251;
// bram[11877] = 253;
// bram[11878] = 253;
// bram[11879] = 252;
// bram[11880] = 248;
// bram[11881] = 244;
// bram[11882] = 237;
// bram[11883] = 229;
// bram[11884] = 220;
// bram[11885] = 209;
// bram[11886] = 198;
// bram[11887] = 185;
// bram[11888] = 172;
// bram[11889] = 158;
// bram[11890] = 143;
// bram[11891] = 129;
// bram[11892] = 114;
// bram[11893] = 100;
// bram[11894] = 86;
// bram[11895] = 72;
// bram[11896] = 59;
// bram[11897] = 47;
// bram[11898] = 36;
// bram[11899] = 27;
// bram[11900] = 18;
// bram[11901] = 11;
// bram[11902] = 6;
// bram[11903] = 2;
// bram[11904] = 0;
// bram[11905] = 0;
// bram[11906] = 1;
// bram[11907] = 4;
// bram[11908] = 8;
// bram[11909] = 14;
// bram[11910] = 22;
// bram[11911] = 31;
// bram[11912] = 41;
// bram[11913] = 53;
// bram[11914] = 65;
// bram[11915] = 78;
// bram[11916] = 92;
// bram[11917] = 107;
// bram[11918] = 121;
// bram[11919] = 136;
// bram[11920] = 150;
// bram[11921] = 165;
// bram[11922] = 178;
// bram[11923] = 191;
// bram[11924] = 203;
// bram[11925] = 215;
// bram[11926] = 224;
// bram[11927] = 233;
// bram[11928] = 240;
// bram[11929] = 246;
// bram[11930] = 250;
// bram[11931] = 253;
// bram[11932] = 253;
// bram[11933] = 253;
// bram[11934] = 250;
// bram[11935] = 246;
// bram[11936] = 240;
// bram[11937] = 233;
// bram[11938] = 224;
// bram[11939] = 214;
// bram[11940] = 203;
// bram[11941] = 191;
// bram[11942] = 177;
// bram[11943] = 164;
// bram[11944] = 150;
// bram[11945] = 135;
// bram[11946] = 120;
// bram[11947] = 106;
// bram[11948] = 91;
// bram[11949] = 78;
// bram[11950] = 64;
// bram[11951] = 52;
// bram[11952] = 41;
// bram[11953] = 31;
// bram[11954] = 22;
// bram[11955] = 14;
// bram[11956] = 8;
// bram[11957] = 4;
// bram[11958] = 1;
// bram[11959] = 0;
// bram[11960] = 0;
// bram[11961] = 2;
// bram[11962] = 6;
// bram[11963] = 12;
// bram[11964] = 19;
// bram[11965] = 27;
// bram[11966] = 37;
// bram[11967] = 48;
// bram[11968] = 60;
// bram[11969] = 73;
// bram[11970] = 86;
// bram[11971] = 100;
// bram[11972] = 115;
// bram[11973] = 130;
// bram[11974] = 144;
// bram[11975] = 159;
// bram[11976] = 173;
// bram[11977] = 186;
// bram[11978] = 198;
// bram[11979] = 210;
// bram[11980] = 220;
// bram[11981] = 230;
// bram[11982] = 238;
// bram[11983] = 244;
// bram[11984] = 249;
// bram[11985] = 252;
// bram[11986] = 253;
// bram[11987] = 253;
// bram[11988] = 251;
// bram[11989] = 248;
// bram[11990] = 243;
// bram[11991] = 236;
// bram[11992] = 228;
// bram[11993] = 218;
// bram[11994] = 208;
// bram[11995] = 196;
// bram[11996] = 183;
// bram[11997] = 170;
// bram[11998] = 156;
// bram[11999] = 141;
// bram[12000] = 126;
// bram[12001] = 112;
// bram[12002] = 97;
// bram[12003] = 83;
// bram[12004] = 70;
// bram[12005] = 57;
// bram[12006] = 45;
// bram[12007] = 35;
// bram[12008] = 25;
// bram[12009] = 17;
// bram[12010] = 10;
// bram[12011] = 5;
// bram[12012] = 2;
// bram[12013] = 0;
// bram[12014] = 0;
// bram[12015] = 1;
// bram[12016] = 4;
// bram[12017] = 9;
// bram[12018] = 15;
// bram[12019] = 23;
// bram[12020] = 33;
// bram[12021] = 43;
// bram[12022] = 55;
// bram[12023] = 67;
// bram[12024] = 80;
// bram[12025] = 94;
// bram[12026] = 109;
// bram[12027] = 123;
// bram[12028] = 138;
// bram[12029] = 153;
// bram[12030] = 167;
// bram[12031] = 180;
// bram[12032] = 193;
// bram[12033] = 205;
// bram[12034] = 216;
// bram[12035] = 226;
// bram[12036] = 234;
// bram[12037] = 241;
// bram[12038] = 247;
// bram[12039] = 251;
// bram[12040] = 253;
// bram[12041] = 253;
// bram[12042] = 252;
// bram[12043] = 249;
// bram[12044] = 245;
// bram[12045] = 239;
// bram[12046] = 231;
// bram[12047] = 222;
// bram[12048] = 212;
// bram[12049] = 201;
// bram[12050] = 189;
// bram[12051] = 175;
// bram[12052] = 162;
// bram[12053] = 147;
// bram[12054] = 133;
// bram[12055] = 118;
// bram[12056] = 103;
// bram[12057] = 89;
// bram[12058] = 76;
// bram[12059] = 62;
// bram[12060] = 50;
// bram[12061] = 39;
// bram[12062] = 29;
// bram[12063] = 20;
// bram[12064] = 13;
// bram[12065] = 7;
// bram[12066] = 3;
// bram[12067] = 0;
// bram[12068] = 0;
// bram[12069] = 0;
// bram[12070] = 3;
// bram[12071] = 7;
// bram[12072] = 13;
// bram[12073] = 20;
// bram[12074] = 29;
// bram[12075] = 38;
// bram[12076] = 50;
// bram[12077] = 62;
// bram[12078] = 75;
// bram[12079] = 88;
// bram[12080] = 103;
// bram[12081] = 117;
// bram[12082] = 132;
// bram[12083] = 146;
// bram[12084] = 161;
// bram[12085] = 175;
// bram[12086] = 188;
// bram[12087] = 200;
// bram[12088] = 212;
// bram[12089] = 222;
// bram[12090] = 231;
// bram[12091] = 239;
// bram[12092] = 245;
// bram[12093] = 249;
// bram[12094] = 252;
// bram[12095] = 253;
// bram[12096] = 253;
// bram[12097] = 251;
// bram[12098] = 247;
// bram[12099] = 242;
// bram[12100] = 235;
// bram[12101] = 226;
// bram[12102] = 217;
// bram[12103] = 206;
// bram[12104] = 194;
// bram[12105] = 181;
// bram[12106] = 167;
// bram[12107] = 153;
// bram[12108] = 139;
// bram[12109] = 124;
// bram[12110] = 110;
// bram[12111] = 95;
// bram[12112] = 81;
// bram[12113] = 68;
// bram[12114] = 55;
// bram[12115] = 44;
// bram[12116] = 33;
// bram[12117] = 24;
// bram[12118] = 16;
// bram[12119] = 9;
// bram[12120] = 5;
// bram[12121] = 1;
// bram[12122] = 0;
// bram[12123] = 0;
// bram[12124] = 2;
// bram[12125] = 5;
// bram[12126] = 10;
// bram[12127] = 17;
// bram[12128] = 25;
// bram[12129] = 34;
// bram[12130] = 45;
// bram[12131] = 57;
// bram[12132] = 69;
// bram[12133] = 83;
// bram[12134] = 97;
// bram[12135] = 111;
// bram[12136] = 126;
// bram[12137] = 140;
// bram[12138] = 155;
// bram[12139] = 169;
// bram[12140] = 182;
// bram[12141] = 195;
// bram[12142] = 207;
// bram[12143] = 218;
// bram[12144] = 227;
// bram[12145] = 236;
// bram[12146] = 242;
// bram[12147] = 248;
// bram[12148] = 251;
// bram[12149] = 253;
// bram[12150] = 253;
// bram[12151] = 252;
// bram[12152] = 249;
// bram[12153] = 244;
// bram[12154] = 238;
// bram[12155] = 230;
// bram[12156] = 221;
// bram[12157] = 211;
// bram[12158] = 199;
// bram[12159] = 187;
// bram[12160] = 173;
// bram[12161] = 159;
// bram[12162] = 145;
// bram[12163] = 130;
// bram[12164] = 116;
// bram[12165] = 101;
// bram[12166] = 87;
// bram[12167] = 73;
// bram[12168] = 60;
// bram[12169] = 48;
// bram[12170] = 37;
// bram[12171] = 28;
// bram[12172] = 19;
// bram[12173] = 12;
// bram[12174] = 6;
// bram[12175] = 2;
// bram[12176] = 0;
// bram[12177] = 0;
// bram[12178] = 1;
// bram[12179] = 3;
// bram[12180] = 8;
// bram[12181] = 14;
// bram[12182] = 21;
// bram[12183] = 30;
// bram[12184] = 40;
// bram[12185] = 51;
// bram[12186] = 64;
// bram[12187] = 77;
// bram[12188] = 91;
// bram[12189] = 105;
// bram[12190] = 120;
// bram[12191] = 134;
// bram[12192] = 149;
// bram[12193] = 163;
// bram[12194] = 177;
// bram[12195] = 190;
// bram[12196] = 202;
// bram[12197] = 213;
// bram[12198] = 223;
// bram[12199] = 232;
// bram[12200] = 240;
// bram[12201] = 246;
// bram[12202] = 250;
// bram[12203] = 253;
// bram[12204] = 253;
// bram[12205] = 253;
// bram[12206] = 250;
// bram[12207] = 246;
// bram[12208] = 241;
// bram[12209] = 234;
// bram[12210] = 225;
// bram[12211] = 215;
// bram[12212] = 204;
// bram[12213] = 192;
// bram[12214] = 179;
// bram[12215] = 165;
// bram[12216] = 151;
// bram[12217] = 137;
// bram[12218] = 122;
// bram[12219] = 107;
// bram[12220] = 93;
// bram[12221] = 79;
// bram[12222] = 66;
// bram[12223] = 53;
// bram[12224] = 42;
// bram[12225] = 32;
// bram[12226] = 22;
// bram[12227] = 15;
// bram[12228] = 9;
// bram[12229] = 4;
// bram[12230] = 1;
// bram[12231] = 0;
// bram[12232] = 0;
// bram[12233] = 2;
// bram[12234] = 6;
// bram[12235] = 11;
// bram[12236] = 18;
// bram[12237] = 26;
// bram[12238] = 36;
// bram[12239] = 47;
// bram[12240] = 58;
// bram[12241] = 71;
// bram[12242] = 85;
// bram[12243] = 99;
// bram[12244] = 113;
// bram[12245] = 128;
// bram[12246] = 143;
// bram[12247] = 157;
// bram[12248] = 171;
// bram[12249] = 184;
// bram[12250] = 197;
// bram[12251] = 209;
// bram[12252] = 219;
// bram[12253] = 229;
// bram[12254] = 237;
// bram[12255] = 243;
// bram[12256] = 248;
// bram[12257] = 252;
// bram[12258] = 253;
// bram[12259] = 253;
// bram[12260] = 252;
// bram[12261] = 248;
// bram[12262] = 243;
// bram[12263] = 237;
// bram[12264] = 229;
// bram[12265] = 219;
// bram[12266] = 209;
// bram[12267] = 197;
// bram[12268] = 185;
// bram[12269] = 171;
// bram[12270] = 157;
// bram[12271] = 143;
// bram[12272] = 128;
// bram[12273] = 113;
// bram[12274] = 99;
// bram[12275] = 85;
// bram[12276] = 71;
// bram[12277] = 59;
// bram[12278] = 47;
// bram[12279] = 36;
// bram[12280] = 26;
// bram[12281] = 18;
// bram[12282] = 11;
// bram[12283] = 6;
// bram[12284] = 2;
// bram[12285] = 0;
// bram[12286] = 0;
// bram[12287] = 1;
// bram[12288] = 4;
// bram[12289] = 9;
// bram[12290] = 15;
// bram[12291] = 22;
// bram[12292] = 32;
// bram[12293] = 42;
// bram[12294] = 53;
// bram[12295] = 66;
// bram[12296] = 79;
// bram[12297] = 93;
// bram[12298] = 107;
// bram[12299] = 122;
// bram[12300] = 136;
// bram[12301] = 151;
// bram[12302] = 165;
// bram[12303] = 179;
// bram[12304] = 192;
// bram[12305] = 204;
// bram[12306] = 215;
// bram[12307] = 225;
// bram[12308] = 234;
// bram[12309] = 241;
// bram[12310] = 246;
// bram[12311] = 250;
// bram[12312] = 253;
// bram[12313] = 253;
// bram[12314] = 253;
// bram[12315] = 250;
// bram[12316] = 246;
// bram[12317] = 240;
// bram[12318] = 232;
// bram[12319] = 224;
// bram[12320] = 213;
// bram[12321] = 202;
// bram[12322] = 190;
// bram[12323] = 177;
// bram[12324] = 163;
// bram[12325] = 149;
// bram[12326] = 134;
// bram[12327] = 120;
// bram[12328] = 105;
// bram[12329] = 91;
// bram[12330] = 77;
// bram[12331] = 64;
// bram[12332] = 52;
// bram[12333] = 40;
// bram[12334] = 30;
// bram[12335] = 21;
// bram[12336] = 14;
// bram[12337] = 8;
// bram[12338] = 3;
// bram[12339] = 1;
// bram[12340] = 0;
// bram[12341] = 0;
// bram[12342] = 2;
// bram[12343] = 6;
// bram[12344] = 12;
// bram[12345] = 19;
// bram[12346] = 28;
// bram[12347] = 37;
// bram[12348] = 48;
// bram[12349] = 60;
// bram[12350] = 73;
// bram[12351] = 87;
// bram[12352] = 101;
// bram[12353] = 116;
// bram[12354] = 130;
// bram[12355] = 145;
// bram[12356] = 159;
// bram[12357] = 173;
// bram[12358] = 186;
// bram[12359] = 199;
// bram[12360] = 210;
// bram[12361] = 221;
// bram[12362] = 230;
// bram[12363] = 238;
// bram[12364] = 244;
// bram[12365] = 249;
// bram[12366] = 252;
// bram[12367] = 253;
// bram[12368] = 253;
// bram[12369] = 251;
// bram[12370] = 248;
// bram[12371] = 242;
// bram[12372] = 236;
// bram[12373] = 227;
// bram[12374] = 218;
// bram[12375] = 207;
// bram[12376] = 195;
// bram[12377] = 182;
// bram[12378] = 169;
// bram[12379] = 155;
// bram[12380] = 140;
// bram[12381] = 126;
// bram[12382] = 111;
// bram[12383] = 97;
// bram[12384] = 83;
// bram[12385] = 69;
// bram[12386] = 57;
// bram[12387] = 45;
// bram[12388] = 34;
// bram[12389] = 25;
// bram[12390] = 17;
// bram[12391] = 10;
// bram[12392] = 5;
// bram[12393] = 2;
// bram[12394] = 0;
// bram[12395] = 0;
// bram[12396] = 1;
// bram[12397] = 5;
// bram[12398] = 9;
// bram[12399] = 16;
// bram[12400] = 24;
// bram[12401] = 33;
// bram[12402] = 44;
// bram[12403] = 55;
// bram[12404] = 68;
// bram[12405] = 81;
// bram[12406] = 95;
// bram[12407] = 109;
// bram[12408] = 124;
// bram[12409] = 139;
// bram[12410] = 153;
// bram[12411] = 167;
// bram[12412] = 181;
// bram[12413] = 194;
// bram[12414] = 206;
// bram[12415] = 217;
// bram[12416] = 226;
// bram[12417] = 235;
// bram[12418] = 242;
// bram[12419] = 247;
// bram[12420] = 251;
// bram[12421] = 253;
// bram[12422] = 253;
// bram[12423] = 252;
// bram[12424] = 249;
// bram[12425] = 245;
// bram[12426] = 239;
// bram[12427] = 231;
// bram[12428] = 222;
// bram[12429] = 212;
// bram[12430] = 200;
// bram[12431] = 188;
// bram[12432] = 175;
// bram[12433] = 161;
// bram[12434] = 147;
// bram[12435] = 132;
// bram[12436] = 117;
// bram[12437] = 103;
// bram[12438] = 89;
// bram[12439] = 75;
// bram[12440] = 62;
// bram[12441] = 50;
// bram[12442] = 39;
// bram[12443] = 29;
// bram[12444] = 20;
// bram[12445] = 13;
// bram[12446] = 7;
// bram[12447] = 3;
// bram[12448] = 0;
// bram[12449] = 0;
// bram[12450] = 0;
// bram[12451] = 3;
// bram[12452] = 7;
// bram[12453] = 13;
// bram[12454] = 20;
// bram[12455] = 29;
// bram[12456] = 39;
// bram[12457] = 50;
// bram[12458] = 62;
// bram[12459] = 75;
// bram[12460] = 89;
// bram[12461] = 103;
// bram[12462] = 118;
// bram[12463] = 133;
// bram[12464] = 147;
// bram[12465] = 161;
// bram[12466] = 175;
// bram[12467] = 188;
// bram[12468] = 201;
// bram[12469] = 212;
// bram[12470] = 222;
// bram[12471] = 231;
// bram[12472] = 239;
// bram[12473] = 245;
// bram[12474] = 249;
// bram[12475] = 252;
// bram[12476] = 253;
// bram[12477] = 253;
// bram[12478] = 251;
// bram[12479] = 247;
// bram[12480] = 241;
// bram[12481] = 234;
// bram[12482] = 226;
// bram[12483] = 216;
// bram[12484] = 205;
// bram[12485] = 193;
// bram[12486] = 180;
// bram[12487] = 167;
// bram[12488] = 153;
// bram[12489] = 138;
// bram[12490] = 124;
// bram[12491] = 109;
// bram[12492] = 95;
// bram[12493] = 81;
// bram[12494] = 67;
// bram[12495] = 55;
// bram[12496] = 43;
// bram[12497] = 33;
// bram[12498] = 23;
// bram[12499] = 16;
// bram[12500] = 9;
// bram[12501] = 4;
// bram[12502] = 1;
// bram[12503] = 0;
// bram[12504] = 0;
// bram[12505] = 2;
// bram[12506] = 5;
// bram[12507] = 10;
// bram[12508] = 17;
// bram[12509] = 25;
// bram[12510] = 35;
// bram[12511] = 45;
// bram[12512] = 57;
// bram[12513] = 70;
// bram[12514] = 83;
// bram[12515] = 97;
// bram[12516] = 112;
// bram[12517] = 126;
// bram[12518] = 141;
// bram[12519] = 155;
// bram[12520] = 170;
// bram[12521] = 183;
// bram[12522] = 196;
// bram[12523] = 208;
// bram[12524] = 218;
// bram[12525] = 228;
// bram[12526] = 236;
// bram[12527] = 243;
// bram[12528] = 248;
// bram[12529] = 251;
// bram[12530] = 253;
// bram[12531] = 253;
// bram[12532] = 252;
// bram[12533] = 249;
// bram[12534] = 244;
// bram[12535] = 238;
// bram[12536] = 230;
// bram[12537] = 221;
// bram[12538] = 210;
// bram[12539] = 198;
// bram[12540] = 186;
// bram[12541] = 173;
// bram[12542] = 159;
// bram[12543] = 144;
// bram[12544] = 130;
// bram[12545] = 115;
// bram[12546] = 101;
// bram[12547] = 86;
// bram[12548] = 73;
// bram[12549] = 60;
// bram[12550] = 48;
// bram[12551] = 37;
// bram[12552] = 27;
// bram[12553] = 19;
// bram[12554] = 12;
// bram[12555] = 6;
// bram[12556] = 2;
// bram[12557] = 0;
// bram[12558] = 0;
// bram[12559] = 1;
// bram[12560] = 3;
// bram[12561] = 8;
// bram[12562] = 14;
// bram[12563] = 22;
// bram[12564] = 30;
// bram[12565] = 41;
// bram[12566] = 52;
// bram[12567] = 64;
// bram[12568] = 78;
// bram[12569] = 91;
// bram[12570] = 106;
// bram[12571] = 120;
// bram[12572] = 135;
// bram[12573] = 149;
// bram[12574] = 164;
// bram[12575] = 177;
// bram[12576] = 190;
// bram[12577] = 203;
// bram[12578] = 214;
// bram[12579] = 224;
// bram[12580] = 233;
// bram[12581] = 240;
// bram[12582] = 246;
// bram[12583] = 250;
// bram[12584] = 253;
// bram[12585] = 253;
// bram[12586] = 253;
// bram[12587] = 250;
// bram[12588] = 246;
// bram[12589] = 240;
// bram[12590] = 233;
// bram[12591] = 225;
// bram[12592] = 215;
// bram[12593] = 203;
// bram[12594] = 191;
// bram[12595] = 178;
// bram[12596] = 165;
// bram[12597] = 150;
// bram[12598] = 136;
// bram[12599] = 121;
// bram[12600] = 107;
// bram[12601] = 92;
// bram[12602] = 78;
// bram[12603] = 65;
// bram[12604] = 53;
// bram[12605] = 41;
// bram[12606] = 31;
// bram[12607] = 22;
// bram[12608] = 14;
// bram[12609] = 8;
// bram[12610] = 4;
// bram[12611] = 1;
// bram[12612] = 0;
// bram[12613] = 0;
// bram[12614] = 2;
// bram[12615] = 6;
// bram[12616] = 11;
// bram[12617] = 18;
// bram[12618] = 27;
// bram[12619] = 36;
// bram[12620] = 47;
// bram[12621] = 59;
// bram[12622] = 72;
// bram[12623] = 85;
// bram[12624] = 100;
// bram[12625] = 114;
// bram[12626] = 129;
// bram[12627] = 143;
// bram[12628] = 158;
// bram[12629] = 172;
// bram[12630] = 185;
// bram[12631] = 198;
// bram[12632] = 209;
// bram[12633] = 220;
// bram[12634] = 229;
// bram[12635] = 237;
// bram[12636] = 244;
// bram[12637] = 248;
// bram[12638] = 252;
// bram[12639] = 253;
// bram[12640] = 253;
// bram[12641] = 251;
// bram[12642] = 248;
// bram[12643] = 243;
// bram[12644] = 236;
// bram[12645] = 228;
// bram[12646] = 219;
// bram[12647] = 208;
// bram[12648] = 197;
// bram[12649] = 184;
// bram[12650] = 170;
// bram[12651] = 156;
// bram[12652] = 142;
// bram[12653] = 127;
// bram[12654] = 113;
// bram[12655] = 98;
// bram[12656] = 84;
// bram[12657] = 71;
// bram[12658] = 58;
// bram[12659] = 46;
// bram[12660] = 35;
// bram[12661] = 26;
// bram[12662] = 17;
// bram[12663] = 11;
// bram[12664] = 5;
// bram[12665] = 2;
// bram[12666] = 0;
// bram[12667] = 0;
// bram[12668] = 1;
// bram[12669] = 4;
// bram[12670] = 9;
// bram[12671] = 15;
// bram[12672] = 23;
// bram[12673] = 32;
// bram[12674] = 42;
// bram[12675] = 54;
// bram[12676] = 66;
// bram[12677] = 80;
// bram[12678] = 94;
// bram[12679] = 108;
// bram[12680] = 123;
// bram[12681] = 137;
// bram[12682] = 152;
// bram[12683] = 166;
// bram[12684] = 179;
// bram[12685] = 192;
// bram[12686] = 204;
// bram[12687] = 216;
// bram[12688] = 225;
// bram[12689] = 234;
// bram[12690] = 241;
// bram[12691] = 247;
// bram[12692] = 251;
// bram[12693] = 253;
// bram[12694] = 253;
// bram[12695] = 252;
// bram[12696] = 250;
// bram[12697] = 245;
// bram[12698] = 239;
// bram[12699] = 232;
// bram[12700] = 223;
// bram[12701] = 213;
// bram[12702] = 202;
// bram[12703] = 189;
// bram[12704] = 176;
// bram[12705] = 162;
// bram[12706] = 148;
// bram[12707] = 134;
// bram[12708] = 119;
// bram[12709] = 104;
// bram[12710] = 90;
// bram[12711] = 76;
// bram[12712] = 63;
// bram[12713] = 51;
// bram[12714] = 40;
// bram[12715] = 30;
// bram[12716] = 21;
// bram[12717] = 13;
// bram[12718] = 7;
// bram[12719] = 3;
// bram[12720] = 1;
// bram[12721] = 0;
// bram[12722] = 0;
// bram[12723] = 3;
// bram[12724] = 7;
// bram[12725] = 12;
// bram[12726] = 19;
// bram[12727] = 28;
// bram[12728] = 38;
// bram[12729] = 49;
// bram[12730] = 61;
// bram[12731] = 74;
// bram[12732] = 88;
// bram[12733] = 102;
// bram[12734] = 116;
// bram[12735] = 131;
// bram[12736] = 146;
// bram[12737] = 160;
// bram[12738] = 174;
// bram[12739] = 187;
// bram[12740] = 200;
// bram[12741] = 211;
// bram[12742] = 221;
// bram[12743] = 230;
// bram[12744] = 238;
// bram[12745] = 244;
// bram[12746] = 249;
// bram[12747] = 252;
// bram[12748] = 253;
// bram[12749] = 253;
// bram[12750] = 251;
// bram[12751] = 247;
// bram[12752] = 242;
// bram[12753] = 235;
// bram[12754] = 227;
// bram[12755] = 217;
// bram[12756] = 207;
// bram[12757] = 195;
// bram[12758] = 182;
// bram[12759] = 168;
// bram[12760] = 154;
// bram[12761] = 140;
// bram[12762] = 125;
// bram[12763] = 110;
// bram[12764] = 96;
// bram[12765] = 82;
// bram[12766] = 69;
// bram[12767] = 56;
// bram[12768] = 44;
// bram[12769] = 34;
// bram[12770] = 24;
// bram[12771] = 16;
// bram[12772] = 10;
// bram[12773] = 5;
// bram[12774] = 1;
// bram[12775] = 0;
// bram[12776] = 0;
// bram[12777] = 1;
// bram[12778] = 5;
// bram[12779] = 10;
// bram[12780] = 16;
// bram[12781] = 24;
// bram[12782] = 34;
// bram[12783] = 44;
// bram[12784] = 56;
// bram[12785] = 68;
// bram[12786] = 82;
// bram[12787] = 96;
// bram[12788] = 110;
// bram[12789] = 125;
// bram[12790] = 139;
// bram[12791] = 154;
// bram[12792] = 168;
// bram[12793] = 182;
// bram[12794] = 194;
// bram[12795] = 206;
// bram[12796] = 217;
// bram[12797] = 227;
// bram[12798] = 235;
// bram[12799] = 242;
// bram[12800] = 247;
// bram[12801] = 251;
// bram[12802] = 253;
// bram[12803] = 253;
// bram[12804] = 252;
// bram[12805] = 249;
// bram[12806] = 245;
// bram[12807] = 238;
// bram[12808] = 231;
// bram[12809] = 222;
// bram[12810] = 211;
// bram[12811] = 200;
// bram[12812] = 187;
// bram[12813] = 174;
// bram[12814] = 160;
// bram[12815] = 146;
// bram[12816] = 131;
// bram[12817] = 117;
// bram[12818] = 102;
// bram[12819] = 88;
// bram[12820] = 74;
// bram[12821] = 61;
// bram[12822] = 49;
// bram[12823] = 38;
// bram[12824] = 28;
// bram[12825] = 20;
// bram[12826] = 12;
// bram[12827] = 7;
// bram[12828] = 3;
// bram[12829] = 0;
// bram[12830] = 0;
// bram[12831] = 0;
// bram[12832] = 3;
// bram[12833] = 7;
// bram[12834] = 13;
// bram[12835] = 21;
// bram[12836] = 29;
// bram[12837] = 39;
// bram[12838] = 51;
// bram[12839] = 63;
// bram[12840] = 76;
// bram[12841] = 90;
// bram[12842] = 104;
// bram[12843] = 119;
// bram[12844] = 133;
// bram[12845] = 148;
// bram[12846] = 162;
// bram[12847] = 176;
// bram[12848] = 189;
// bram[12849] = 201;
// bram[12850] = 213;
// bram[12851] = 223;
// bram[12852] = 232;
// bram[12853] = 239;
// bram[12854] = 245;
// bram[12855] = 250;
// bram[12856] = 252;
// bram[12857] = 253;
// bram[12858] = 253;
// bram[12859] = 251;
// bram[12860] = 247;
// bram[12861] = 241;
// bram[12862] = 234;
// bram[12863] = 226;
// bram[12864] = 216;
// bram[12865] = 205;
// bram[12866] = 193;
// bram[12867] = 180;
// bram[12868] = 166;
// bram[12869] = 152;
// bram[12870] = 137;
// bram[12871] = 123;
// bram[12872] = 108;
// bram[12873] = 94;
// bram[12874] = 80;
// bram[12875] = 67;
// bram[12876] = 54;
// bram[12877] = 43;
// bram[12878] = 32;
// bram[12879] = 23;
// bram[12880] = 15;
// bram[12881] = 9;
// bram[12882] = 4;
// bram[12883] = 1;
// bram[12884] = 0;
// bram[12885] = 0;
// bram[12886] = 2;
// bram[12887] = 5;
// bram[12888] = 11;
// bram[12889] = 17;
// bram[12890] = 26;
// bram[12891] = 35;
// bram[12892] = 46;
// bram[12893] = 58;
// bram[12894] = 70;
// bram[12895] = 84;
// bram[12896] = 98;
// bram[12897] = 112;
// bram[12898] = 127;
// bram[12899] = 142;
// bram[12900] = 156;
// bram[12901] = 170;
// bram[12902] = 184;
// bram[12903] = 196;
// bram[12904] = 208;
// bram[12905] = 219;
// bram[12906] = 228;
// bram[12907] = 236;
// bram[12908] = 243;
// bram[12909] = 248;
// bram[12910] = 251;
// bram[12911] = 253;
// bram[12912] = 253;
// bram[12913] = 252;
// bram[12914] = 249;
// bram[12915] = 244;
// bram[12916] = 237;
// bram[12917] = 229;
// bram[12918] = 220;
// bram[12919] = 210;
// bram[12920] = 198;
// bram[12921] = 185;
// bram[12922] = 172;
// bram[12923] = 158;
// bram[12924] = 144;
// bram[12925] = 129;
// bram[12926] = 114;
// bram[12927] = 100;
// bram[12928] = 86;
// bram[12929] = 72;
// bram[12930] = 59;
// bram[12931] = 47;
// bram[12932] = 36;
// bram[12933] = 27;
// bram[12934] = 18;
// bram[12935] = 11;
// bram[12936] = 6;
// bram[12937] = 2;
// bram[12938] = 0;
// bram[12939] = 0;
// bram[12940] = 1;
// bram[12941] = 4;
// bram[12942] = 8;
// bram[12943] = 14;
// bram[12944] = 22;
// bram[12945] = 31;
// bram[12946] = 41;
// bram[12947] = 53;
// bram[12948] = 65;
// bram[12949] = 78;
// bram[12950] = 92;
// bram[12951] = 106;
// bram[12952] = 121;
// bram[12953] = 136;
// bram[12954] = 150;
// bram[12955] = 164;
// bram[12956] = 178;
// bram[12957] = 191;
// bram[12958] = 203;
// bram[12959] = 214;
// bram[12960] = 224;
// bram[12961] = 233;
// bram[12962] = 240;
// bram[12963] = 246;
// bram[12964] = 250;
// bram[12965] = 253;
// bram[12966] = 253;
// bram[12967] = 253;
// bram[12968] = 250;
// bram[12969] = 246;
// bram[12970] = 240;
// bram[12971] = 233;
// bram[12972] = 224;
// bram[12973] = 214;
// bram[12974] = 203;
// bram[12975] = 191;
// bram[12976] = 178;
// bram[12977] = 164;
// bram[12978] = 150;
// bram[12979] = 135;
// bram[12980] = 121;
// bram[12981] = 106;
// bram[12982] = 92;
// bram[12983] = 78;
// bram[12984] = 65;
// bram[12985] = 52;
// bram[12986] = 41;
// bram[12987] = 31;
// bram[12988] = 22;
// bram[12989] = 14;
// bram[12990] = 8;
// bram[12991] = 4;
// bram[12992] = 1;
// bram[12993] = 0;
// bram[12994] = 0;
// bram[12995] = 2;
// bram[12996] = 6;
// bram[12997] = 12;
// bram[12998] = 19;
// bram[12999] = 27;
// bram[13000] = 37;
// bram[13001] = 48;
// bram[13002] = 60;
// bram[13003] = 73;
// bram[13004] = 86;
// bram[13005] = 100;
// bram[13006] = 115;
// bram[13007] = 129;
// bram[13008] = 144;
// bram[13009] = 158;
// bram[13010] = 172;
// bram[13011] = 186;
// bram[13012] = 198;
// bram[13013] = 210;
// bram[13014] = 220;
// bram[13015] = 230;
// bram[13016] = 237;
// bram[13017] = 244;
// bram[13018] = 249;
// bram[13019] = 252;
// bram[13020] = 253;
// bram[13021] = 253;
// bram[13022] = 251;
// bram[13023] = 248;
// bram[13024] = 243;
// bram[13025] = 236;
// bram[13026] = 228;
// bram[13027] = 218;
// bram[13028] = 208;
// bram[13029] = 196;
// bram[13030] = 183;
// bram[13031] = 170;
// bram[13032] = 156;
// bram[13033] = 141;
// bram[13034] = 127;
// bram[13035] = 112;
// bram[13036] = 98;
// bram[13037] = 84;
// bram[13038] = 70;
// bram[13039] = 57;
// bram[13040] = 46;
// bram[13041] = 35;
// bram[13042] = 25;
// bram[13043] = 17;
// bram[13044] = 10;
// bram[13045] = 5;
// bram[13046] = 2;
// bram[13047] = 0;
// bram[13048] = 0;
// bram[13049] = 1;
// bram[13050] = 4;
// bram[13051] = 9;
// bram[13052] = 15;
// bram[13053] = 23;
// bram[13054] = 32;
// bram[13055] = 43;
// bram[13056] = 54;
// bram[13057] = 67;
// bram[13058] = 80;
// bram[13059] = 94;
// bram[13060] = 109;
// bram[13061] = 123;
// bram[13062] = 138;
// bram[13063] = 152;
// bram[13064] = 167;
// bram[13065] = 180;
// bram[13066] = 193;
// bram[13067] = 205;
// bram[13068] = 216;
// bram[13069] = 226;
// bram[13070] = 234;
// bram[13071] = 241;
// bram[13072] = 247;
// bram[13073] = 251;
// bram[13074] = 253;
// bram[13075] = 253;
// bram[13076] = 252;
// bram[13077] = 250;
// bram[13078] = 245;
// bram[13079] = 239;
// bram[13080] = 232;
// bram[13081] = 223;
// bram[13082] = 212;
// bram[13083] = 201;
// bram[13084] = 189;
// bram[13085] = 176;
// bram[13086] = 162;
// bram[13087] = 147;
// bram[13088] = 133;
// bram[13089] = 118;
// bram[13090] = 104;
// bram[13091] = 89;
// bram[13092] = 76;
// bram[13093] = 63;
// bram[13094] = 50;
// bram[13095] = 39;
// bram[13096] = 29;
// bram[13097] = 20;
// bram[13098] = 13;
// bram[13099] = 7;
// bram[13100] = 3;
// bram[13101] = 0;
// bram[13102] = 0;
// bram[13103] = 0;
// bram[13104] = 3;
// bram[13105] = 7;
// bram[13106] = 13;
// bram[13107] = 20;
// bram[13108] = 28;
// bram[13109] = 38;
// bram[13110] = 49;
// bram[13111] = 62;
// bram[13112] = 75;
// bram[13113] = 88;
// bram[13114] = 103;
// bram[13115] = 117;
// bram[13116] = 132;
// bram[13117] = 146;
// bram[13118] = 161;
// bram[13119] = 174;
// bram[13120] = 188;
// bram[13121] = 200;
// bram[13122] = 212;
// bram[13123] = 222;
// bram[13124] = 231;
// bram[13125] = 239;
// bram[13126] = 245;
// bram[13127] = 249;
// bram[13128] = 252;
// bram[13129] = 253;
// bram[13130] = 253;
// bram[13131] = 251;
// bram[13132] = 247;
// bram[13133] = 242;
// bram[13134] = 235;
// bram[13135] = 227;
// bram[13136] = 217;
// bram[13137] = 206;
// bram[13138] = 194;
// bram[13139] = 181;
// bram[13140] = 168;
// bram[13141] = 154;
// bram[13142] = 139;
// bram[13143] = 124;
// bram[13144] = 110;
// bram[13145] = 95;
// bram[13146] = 81;
// bram[13147] = 68;
// bram[13148] = 55;
// bram[13149] = 44;
// bram[13150] = 33;
// bram[13151] = 24;
// bram[13152] = 16;
// bram[13153] = 10;
// bram[13154] = 5;
// bram[13155] = 1;
// bram[13156] = 0;
// bram[13157] = 0;
// bram[13158] = 1;
// bram[13159] = 5;
// bram[13160] = 10;
// bram[13161] = 17;
// bram[13162] = 25;
// bram[13163] = 34;
// bram[13164] = 45;
// bram[13165] = 56;
// bram[13166] = 69;
// bram[13167] = 82;
// bram[13168] = 96;
// bram[13169] = 111;
// bram[13170] = 126;
// bram[13171] = 140;
// bram[13172] = 155;
// bram[13173] = 169;
// bram[13174] = 182;
// bram[13175] = 195;
// bram[13176] = 207;
// bram[13177] = 218;
// bram[13178] = 227;
// bram[13179] = 235;
// bram[13180] = 242;
// bram[13181] = 247;
// bram[13182] = 251;
// bram[13183] = 253;
// bram[13184] = 253;
// bram[13185] = 252;
// bram[13186] = 249;
// bram[13187] = 244;
// bram[13188] = 238;
// bram[13189] = 230;
// bram[13190] = 221;
// bram[13191] = 211;
// bram[13192] = 199;
// bram[13193] = 187;
// bram[13194] = 173;
// bram[13195] = 160;
// bram[13196] = 145;
// bram[13197] = 131;
// bram[13198] = 116;
// bram[13199] = 101;
// bram[13200] = 87;
// bram[13201] = 74;
// bram[13202] = 61;
// bram[13203] = 49;
// bram[13204] = 38;
// bram[13205] = 28;
// bram[13206] = 19;
// bram[13207] = 12;
// bram[13208] = 6;
// bram[13209] = 2;
// bram[13210] = 0;
// bram[13211] = 0;
// bram[13212] = 1;
// bram[13213] = 3;
// bram[13214] = 8;
// bram[13215] = 14;
// bram[13216] = 21;
// bram[13217] = 30;
// bram[13218] = 40;
// bram[13219] = 51;
// bram[13220] = 64;
// bram[13221] = 77;
// bram[13222] = 90;
// bram[13223] = 105;
// bram[13224] = 119;
// bram[13225] = 134;
// bram[13226] = 149;
// bram[13227] = 163;
// bram[13228] = 177;
// bram[13229] = 190;
// bram[13230] = 202;
// bram[13231] = 213;
// bram[13232] = 223;
// bram[13233] = 232;
// bram[13234] = 240;
// bram[13235] = 245;
// bram[13236] = 250;
// bram[13237] = 252;
// bram[13238] = 253;
// bram[13239] = 253;
// bram[13240] = 250;
// bram[13241] = 246;
// bram[13242] = 241;
// bram[13243] = 234;
// bram[13244] = 225;
// bram[13245] = 215;
// bram[13246] = 204;
// bram[13247] = 192;
// bram[13248] = 179;
// bram[13249] = 165;
// bram[13250] = 151;
// bram[13251] = 137;
// bram[13252] = 122;
// bram[13253] = 108;
// bram[13254] = 93;
// bram[13255] = 79;
// bram[13256] = 66;
// bram[13257] = 54;
// bram[13258] = 42;
// bram[13259] = 32;
// bram[13260] = 23;
// bram[13261] = 15;
// bram[13262] = 9;
// bram[13263] = 4;
// bram[13264] = 1;
// bram[13265] = 0;
// bram[13266] = 0;
// bram[13267] = 2;
// bram[13268] = 6;
// bram[13269] = 11;
// bram[13270] = 18;
// bram[13271] = 26;
// bram[13272] = 36;
// bram[13273] = 46;
// bram[13274] = 58;
// bram[13275] = 71;
// bram[13276] = 85;
// bram[13277] = 99;
// bram[13278] = 113;
// bram[13279] = 128;
// bram[13280] = 142;
// bram[13281] = 157;
// bram[13282] = 171;
// bram[13283] = 184;
// bram[13284] = 197;
// bram[13285] = 209;
// bram[13286] = 219;
// bram[13287] = 229;
// bram[13288] = 237;
// bram[13289] = 243;
// bram[13290] = 248;
// bram[13291] = 252;
// bram[13292] = 253;
// bram[13293] = 253;
// bram[13294] = 252;
// bram[13295] = 248;
// bram[13296] = 243;
// bram[13297] = 237;
// bram[13298] = 229;
// bram[13299] = 220;
// bram[13300] = 209;
// bram[13301] = 197;
// bram[13302] = 185;
// bram[13303] = 171;
// bram[13304] = 157;
// bram[13305] = 143;
// bram[13306] = 128;
// bram[13307] = 114;
// bram[13308] = 99;
// bram[13309] = 85;
// bram[13310] = 72;
// bram[13311] = 59;
// bram[13312] = 47;
// bram[13313] = 36;
// bram[13314] = 26;
// bram[13315] = 18;
// bram[13316] = 11;
// bram[13317] = 6;
// bram[13318] = 2;
// bram[13319] = 0;
// bram[13320] = 0;
// bram[13321] = 1;
// bram[13322] = 4;
// bram[13323] = 8;
// bram[13324] = 15;
// bram[13325] = 22;
// bram[13326] = 31;
// bram[13327] = 42;
// bram[13328] = 53;
// bram[13329] = 66;
// bram[13330] = 79;
// bram[13331] = 93;
// bram[13332] = 107;
// bram[13333] = 122;
// bram[13334] = 136;
// bram[13335] = 151;
// bram[13336] = 165;
// bram[13337] = 179;
// bram[13338] = 192;
// bram[13339] = 204;
// bram[13340] = 215;
// bram[13341] = 225;
// bram[13342] = 233;
// bram[13343] = 241;
// bram[13344] = 246;
// bram[13345] = 250;
// bram[13346] = 253;
// bram[13347] = 253;
// bram[13348] = 253;
// bram[13349] = 250;
// bram[13350] = 246;
// bram[13351] = 240;
// bram[13352] = 232;
// bram[13353] = 224;
// bram[13354] = 214;
// bram[13355] = 202;
// bram[13356] = 190;
// bram[13357] = 177;
// bram[13358] = 163;
// bram[13359] = 149;
// bram[13360] = 134;
// bram[13361] = 120;
// bram[13362] = 105;
// bram[13363] = 91;
// bram[13364] = 77;
// bram[13365] = 64;
// bram[13366] = 52;
// bram[13367] = 40;
// bram[13368] = 30;
// bram[13369] = 21;
// bram[13370] = 14;
// bram[13371] = 8;
// bram[13372] = 3;
// bram[13373] = 1;
// bram[13374] = 0;
// bram[13375] = 0;
// bram[13376] = 2;
// bram[13377] = 6;
// bram[13378] = 12;
// bram[13379] = 19;
// bram[13380] = 27;
// bram[13381] = 37;
// bram[13382] = 48;
// bram[13383] = 60;
// bram[13384] = 73;
// bram[13385] = 87;
// bram[13386] = 101;
// bram[13387] = 115;
// bram[13388] = 130;
// bram[13389] = 145;
// bram[13390] = 159;
// bram[13391] = 173;
// bram[13392] = 186;
// bram[13393] = 199;
// bram[13394] = 210;
// bram[13395] = 221;
// bram[13396] = 230;
// bram[13397] = 238;
// bram[13398] = 244;
// bram[13399] = 249;
// bram[13400] = 252;
// bram[13401] = 253;
// bram[13402] = 253;
// bram[13403] = 251;
// bram[13404] = 248;
// bram[13405] = 242;
// bram[13406] = 236;
// bram[13407] = 228;
// bram[13408] = 218;
// bram[13409] = 207;
// bram[13410] = 195;
// bram[13411] = 183;
// bram[13412] = 169;
// bram[13413] = 155;
// bram[13414] = 141;
// bram[13415] = 126;
// bram[13416] = 111;
// bram[13417] = 97;
// bram[13418] = 83;
// bram[13419] = 69;
// bram[13420] = 57;
// bram[13421] = 45;
// bram[13422] = 34;
// bram[13423] = 25;
// bram[13424] = 17;
// bram[13425] = 10;
// bram[13426] = 5;
// bram[13427] = 2;
// bram[13428] = 0;
// bram[13429] = 0;
// bram[13430] = 1;
// bram[13431] = 4;
// bram[13432] = 9;
// bram[13433] = 16;
// bram[13434] = 24;
// bram[13435] = 33;
// bram[13436] = 43;
// bram[13437] = 55;
// bram[13438] = 68;
// bram[13439] = 81;
// bram[13440] = 95;
// bram[13441] = 109;
// bram[13442] = 124;
// bram[13443] = 139;
// bram[13444] = 153;
// bram[13445] = 167;
// bram[13446] = 181;
// bram[13447] = 194;
// bram[13448] = 206;
// bram[13449] = 217;
// bram[13450] = 226;
// bram[13451] = 235;
// bram[13452] = 242;
// bram[13453] = 247;
// bram[13454] = 251;
// bram[13455] = 253;
// bram[13456] = 253;
// bram[13457] = 252;
// bram[13458] = 249;
// bram[13459] = 245;
// bram[13460] = 239;
// bram[13461] = 231;
// bram[13462] = 222;
// bram[13463] = 212;
// bram[13464] = 201;
// bram[13465] = 188;
// bram[13466] = 175;
// bram[13467] = 161;
// bram[13468] = 147;
// bram[13469] = 132;
// bram[13470] = 118;
// bram[13471] = 103;
// bram[13472] = 89;
// bram[13473] = 75;
// bram[13474] = 62;
// bram[13475] = 50;
// bram[13476] = 39;
// bram[13477] = 29;
// bram[13478] = 20;
// bram[13479] = 13;
// bram[13480] = 7;
// bram[13481] = 3;
// bram[13482] = 0;
// bram[13483] = 0;
// bram[13484] = 0;
// bram[13485] = 3;
// bram[13486] = 7;
// bram[13487] = 13;
// bram[13488] = 20;
// bram[13489] = 29;
// bram[13490] = 39;
// bram[13491] = 50;
// bram[13492] = 62;
// bram[13493] = 75;
// bram[13494] = 89;
// bram[13495] = 103;
// bram[13496] = 118;
// bram[13497] = 132;
// bram[13498] = 147;
// bram[13499] = 161;
// bram[13500] = 175;
// bram[13501] = 188;
// bram[13502] = 201;
// bram[13503] = 212;
// bram[13504] = 222;
// bram[13505] = 231;
// bram[13506] = 239;
// bram[13507] = 245;
// bram[13508] = 249;
// bram[13509] = 252;
// bram[13510] = 253;
// bram[13511] = 253;
// bram[13512] = 251;
// bram[13513] = 247;
// bram[13514] = 241;
// bram[13515] = 235;
// bram[13516] = 226;
// bram[13517] = 216;
// bram[13518] = 205;
// bram[13519] = 193;
// bram[13520] = 181;
// bram[13521] = 167;
// bram[13522] = 153;
// bram[13523] = 138;
// bram[13524] = 124;
// bram[13525] = 109;
// bram[13526] = 95;
// bram[13527] = 81;
// bram[13528] = 67;
// bram[13529] = 55;
// bram[13530] = 43;
// bram[13531] = 33;
// bram[13532] = 24;
// bram[13533] = 16;
// bram[13534] = 9;
// bram[13535] = 4;
// bram[13536] = 1;
// bram[13537] = 0;
// bram[13538] = 0;
// bram[13539] = 2;
// bram[13540] = 5;
// bram[13541] = 10;
// bram[13542] = 17;
// bram[13543] = 25;
// bram[13544] = 34;
// bram[13545] = 45;
// bram[13546] = 57;
// bram[13547] = 70;
// bram[13548] = 83;
// bram[13549] = 97;
// bram[13550] = 112;
// bram[13551] = 126;
// bram[13552] = 141;
// bram[13553] = 155;
// bram[13554] = 169;
// bram[13555] = 183;
// bram[13556] = 196;
// bram[13557] = 207;
// bram[13558] = 218;
// bram[13559] = 228;
// bram[13560] = 236;
// bram[13561] = 243;
// bram[13562] = 248;
// bram[13563] = 251;
// bram[13564] = 253;
// bram[13565] = 253;
// bram[13566] = 252;
// bram[13567] = 249;
// bram[13568] = 244;
// bram[13569] = 238;
// bram[13570] = 230;
// bram[13571] = 221;
// bram[13572] = 210;
// bram[13573] = 199;
// bram[13574] = 186;
// bram[13575] = 173;
// bram[13576] = 159;
// bram[13577] = 144;
// bram[13578] = 130;
// bram[13579] = 115;
// bram[13580] = 101;
// bram[13581] = 87;
// bram[13582] = 73;
// bram[13583] = 60;
// bram[13584] = 48;
// bram[13585] = 37;
// bram[13586] = 27;
// bram[13587] = 19;
// bram[13588] = 12;
// bram[13589] = 6;
// bram[13590] = 2;
// bram[13591] = 0;
// bram[13592] = 0;
// bram[13593] = 1;
// bram[13594] = 3;
// bram[13595] = 8;
// bram[13596] = 14;
// bram[13597] = 21;
// bram[13598] = 30;
// bram[13599] = 41;
// bram[13600] = 52;
// bram[13601] = 64;
// bram[13602] = 77;
// bram[13603] = 91;
// bram[13604] = 105;
// bram[13605] = 120;
// bram[13606] = 135;
// bram[13607] = 149;
// bram[13608] = 163;
// bram[13609] = 177;
// bram[13610] = 190;
// bram[13611] = 203;
// bram[13612] = 214;
// bram[13613] = 224;
// bram[13614] = 233;
// bram[13615] = 240;
// bram[13616] = 246;
// bram[13617] = 250;
// bram[13618] = 253;
// bram[13619] = 253;
// bram[13620] = 253;
// bram[13621] = 250;
// bram[13622] = 246;
// bram[13623] = 241;
// bram[13624] = 233;
// bram[13625] = 225;
// bram[13626] = 215;
// bram[13627] = 204;
// bram[13628] = 191;
// bram[13629] = 178;
// bram[13630] = 165;
// bram[13631] = 151;
// bram[13632] = 136;
// bram[13633] = 121;
// bram[13634] = 107;
// bram[13635] = 93;
// bram[13636] = 79;
// bram[13637] = 65;
// bram[13638] = 53;
// bram[13639] = 42;
// bram[13640] = 31;
// bram[13641] = 22;
// bram[13642] = 15;
// bram[13643] = 8;
// bram[13644] = 4;
// bram[13645] = 1;
// bram[13646] = 0;
// bram[13647] = 0;
// bram[13648] = 2;
// bram[13649] = 6;
// bram[13650] = 11;
// bram[13651] = 18;
// bram[13652] = 26;
// bram[13653] = 36;
// bram[13654] = 47;
// bram[13655] = 59;
// bram[13656] = 72;
// bram[13657] = 85;
// bram[13658] = 99;
// bram[13659] = 114;
// bram[13660] = 128;
// bram[13661] = 143;
// bram[13662] = 158;
// bram[13663] = 171;
// bram[13664] = 185;
// bram[13665] = 197;
// bram[13666] = 209;
// bram[13667] = 220;
// bram[13668] = 229;
// bram[13669] = 237;
// bram[13670] = 243;
// bram[13671] = 248;
// bram[13672] = 252;
// bram[13673] = 253;
// bram[13674] = 253;
// bram[13675] = 252;
// bram[13676] = 248;
// bram[13677] = 243;
// bram[13678] = 237;
// bram[13679] = 228;
// bram[13680] = 219;
// bram[13681] = 208;
// bram[13682] = 197;
// bram[13683] = 184;
// bram[13684] = 171;
// bram[13685] = 157;
// bram[13686] = 142;
// bram[13687] = 128;
// bram[13688] = 113;
// bram[13689] = 99;
// bram[13690] = 84;
// bram[13691] = 71;
// bram[13692] = 58;
// bram[13693] = 46;
// bram[13694] = 35;
// bram[13695] = 26;
// bram[13696] = 18;
// bram[13697] = 11;
// bram[13698] = 6;
// bram[13699] = 2;
// bram[13700] = 0;
// bram[13701] = 0;
// bram[13702] = 1;
// bram[13703] = 4;
// bram[13704] = 9;
// bram[13705] = 15;
// bram[13706] = 23;
// bram[13707] = 32;
// bram[13708] = 42;
// bram[13709] = 54;
// bram[13710] = 66;
// bram[13711] = 79;
// bram[13712] = 93;
// bram[13713] = 108;
// bram[13714] = 122;
// bram[13715] = 137;
// bram[13716] = 151;
// bram[13717] = 166;
// bram[13718] = 179;
// bram[13719] = 192;
// bram[13720] = 204;
// bram[13721] = 215;
// bram[13722] = 225;
// bram[13723] = 234;
// bram[13724] = 241;
// bram[13725] = 246;
// bram[13726] = 250;
// bram[13727] = 253;
// bram[13728] = 253;
// bram[13729] = 252;
// bram[13730] = 250;
// bram[13731] = 245;
// bram[13732] = 239;
// bram[13733] = 232;
// bram[13734] = 223;
// bram[13735] = 213;
// bram[13736] = 202;
// bram[13737] = 190;
// bram[13738] = 176;
// bram[13739] = 163;
// bram[13740] = 148;
// bram[13741] = 134;
// bram[13742] = 119;
// bram[13743] = 105;
// bram[13744] = 90;
// bram[13745] = 77;
// bram[13746] = 63;
// bram[13747] = 51;
// bram[13748] = 40;
// bram[13749] = 30;
// bram[13750] = 21;
// bram[13751] = 13;
// bram[13752] = 8;
// bram[13753] = 3;
// bram[13754] = 1;
// bram[13755] = 0;
// bram[13756] = 0;
// bram[13757] = 3;
// bram[13758] = 7;
// bram[13759] = 12;
// bram[13760] = 19;
// bram[13761] = 28;
// bram[13762] = 38;
// bram[13763] = 49;
// bram[13764] = 61;
// bram[13765] = 74;
// bram[13766] = 87;
// bram[13767] = 102;
// bram[13768] = 116;
// bram[13769] = 131;
// bram[13770] = 145;
// bram[13771] = 160;
// bram[13772] = 174;
// bram[13773] = 187;
// bram[13774] = 199;
// bram[13775] = 211;
// bram[13776] = 221;
// bram[13777] = 230;
// bram[13778] = 238;
// bram[13779] = 244;
// bram[13780] = 249;
// bram[13781] = 252;
// bram[13782] = 253;
// bram[13783] = 253;
// bram[13784] = 251;
// bram[13785] = 247;
// bram[13786] = 242;
// bram[13787] = 235;
// bram[13788] = 227;
// bram[13789] = 217;
// bram[13790] = 207;
// bram[13791] = 195;
// bram[13792] = 182;
// bram[13793] = 168;
// bram[13794] = 154;
// bram[13795] = 140;
// bram[13796] = 125;
// bram[13797] = 111;
// bram[13798] = 96;
// bram[13799] = 82;
// bram[13800] = 69;
// bram[13801] = 56;
// bram[13802] = 44;
// bram[13803] = 34;
// bram[13804] = 24;
// bram[13805] = 16;
// bram[13806] = 10;
// bram[13807] = 5;
// bram[13808] = 1;
// bram[13809] = 0;
// bram[13810] = 0;
// bram[13811] = 1;
// bram[13812] = 5;
// bram[13813] = 10;
// bram[13814] = 16;
// bram[13815] = 24;
// bram[13816] = 33;
// bram[13817] = 44;
// bram[13818] = 56;
// bram[13819] = 68;
// bram[13820] = 82;
// bram[13821] = 96;
// bram[13822] = 110;
// bram[13823] = 125;
// bram[13824] = 139;
// bram[13825] = 154;
// bram[13826] = 168;
// bram[13827] = 181;
// bram[13828] = 194;
// bram[13829] = 206;
// bram[13830] = 217;
// bram[13831] = 227;
// bram[13832] = 235;
// bram[13833] = 242;
// bram[13834] = 247;
// bram[13835] = 251;
// bram[13836] = 253;
// bram[13837] = 253;
// bram[13838] = 252;
// bram[13839] = 249;
// bram[13840] = 245;
// bram[13841] = 238;
// bram[13842] = 231;
// bram[13843] = 222;
// bram[13844] = 211;
// bram[13845] = 200;
// bram[13846] = 188;
// bram[13847] = 174;
// bram[13848] = 160;
// bram[13849] = 146;
// bram[13850] = 131;
// bram[13851] = 117;
// bram[13852] = 102;
// bram[13853] = 88;
// bram[13854] = 74;
// bram[13855] = 61;
// bram[13856] = 49;
// bram[13857] = 38;
// bram[13858] = 28;
// bram[13859] = 20;
// bram[13860] = 12;
// bram[13861] = 7;
// bram[13862] = 3;
// bram[13863] = 0;
// bram[13864] = 0;
// bram[13865] = 0;
// bram[13866] = 3;
// bram[13867] = 7;
// bram[13868] = 13;
// bram[13869] = 21;
// bram[13870] = 29;
// bram[13871] = 39;
// bram[13872] = 51;
// bram[13873] = 63;
// bram[13874] = 76;
// bram[13875] = 90;
// bram[13876] = 104;
// bram[13877] = 118;
// bram[13878] = 133;
// bram[13879] = 148;
// bram[13880] = 162;
// bram[13881] = 176;
// bram[13882] = 189;
// bram[13883] = 201;
// bram[13884] = 213;
// bram[13885] = 223;
// bram[13886] = 232;
// bram[13887] = 239;
// bram[13888] = 245;
// bram[13889] = 250;
// bram[13890] = 252;
// bram[13891] = 253;
// bram[13892] = 253;
// bram[13893] = 251;
// bram[13894] = 247;
// bram[13895] = 241;
// bram[13896] = 234;
// bram[13897] = 226;
// bram[13898] = 216;
// bram[13899] = 205;
// bram[13900] = 193;
// bram[13901] = 180;
// bram[13902] = 166;
// bram[13903] = 152;
// bram[13904] = 138;
// bram[13905] = 123;
// bram[13906] = 108;
// bram[13907] = 94;
// bram[13908] = 80;
// bram[13909] = 67;
// bram[13910] = 54;
// bram[13911] = 43;
// bram[13912] = 32;
// bram[13913] = 23;
// bram[13914] = 15;
// bram[13915] = 9;
// bram[13916] = 4;
// bram[13917] = 1;
// bram[13918] = 0;
// bram[13919] = 0;
// bram[13920] = 2;
// bram[13921] = 5;
// bram[13922] = 11;
// bram[13923] = 17;
// bram[13924] = 25;
// bram[13925] = 35;
// bram[13926] = 46;
// bram[13927] = 58;
// bram[13928] = 70;
// bram[13929] = 84;
// bram[13930] = 98;
// bram[13931] = 112;
// bram[13932] = 127;
// bram[13933] = 142;
// bram[13934] = 156;
// bram[13935] = 170;
// bram[13936] = 183;
// bram[13937] = 196;
// bram[13938] = 208;
// bram[13939] = 219;
// bram[13940] = 228;
// bram[13941] = 236;
// bram[13942] = 243;
// bram[13943] = 248;
// bram[13944] = 251;
// bram[13945] = 253;
// bram[13946] = 253;
// bram[13947] = 252;
// bram[13948] = 249;
// bram[13949] = 244;
// bram[13950] = 237;
// bram[13951] = 229;
// bram[13952] = 220;
// bram[13953] = 210;
// bram[13954] = 198;
// bram[13955] = 185;
// bram[13956] = 172;
// bram[13957] = 158;
// bram[13958] = 144;
// bram[13959] = 129;
// bram[13960] = 115;
// bram[13961] = 100;
// bram[13962] = 86;
// bram[13963] = 72;
// bram[13964] = 59;
// bram[13965] = 47;
// bram[13966] = 37;
// bram[13967] = 27;
// bram[13968] = 18;
// bram[13969] = 11;
// bram[13970] = 6;
// bram[13971] = 2;
// bram[13972] = 0;
// bram[13973] = 0;
// bram[13974] = 1;
// bram[13975] = 4;
// bram[13976] = 8;
// bram[13977] = 14;
// bram[13978] = 22;
// bram[13979] = 31;
// bram[13980] = 41;
// bram[13981] = 52;
// bram[13982] = 65;
// bram[13983] = 78;
// bram[13984] = 92;
// bram[13985] = 106;
// bram[13986] = 121;
// bram[13987] = 135;
// bram[13988] = 150;
// bram[13989] = 164;
// bram[13990] = 178;
// bram[13991] = 191;
// bram[13992] = 203;
// bram[13993] = 214;
// bram[13994] = 224;
// bram[13995] = 233;
// bram[13996] = 240;
// bram[13997] = 246;
// bram[13998] = 250;
// bram[13999] = 253;
// bram[14000] = 254;
// bram[14001] = 253;
// bram[14002] = 250;
// bram[14003] = 246;
// bram[14004] = 240;
// bram[14005] = 233;
// bram[14006] = 224;
// bram[14007] = 214;
// bram[14008] = 203;
// bram[14009] = 191;
// bram[14010] = 178;
// bram[14011] = 164;
// bram[14012] = 150;
// bram[14013] = 135;
// bram[14014] = 121;
// bram[14015] = 106;
// bram[14016] = 92;
// bram[14017] = 78;
// bram[14018] = 65;
// bram[14019] = 52;
// bram[14020] = 41;
// bram[14021] = 31;
// bram[14022] = 22;
// bram[14023] = 14;
// bram[14024] = 8;
// bram[14025] = 4;
// bram[14026] = 1;
// bram[14027] = 0;
// bram[14028] = 0;
// bram[14029] = 2;
// bram[14030] = 6;
// bram[14031] = 11;
// bram[14032] = 18;
// bram[14033] = 27;
// bram[14034] = 37;
// bram[14035] = 47;
// bram[14036] = 59;
// bram[14037] = 72;
// bram[14038] = 86;
// bram[14039] = 100;
// bram[14040] = 115;
// bram[14041] = 129;
// bram[14042] = 144;
// bram[14043] = 158;
// bram[14044] = 172;
// bram[14045] = 185;
// bram[14046] = 198;
// bram[14047] = 210;
// bram[14048] = 220;
// bram[14049] = 229;
// bram[14050] = 237;
// bram[14051] = 244;
// bram[14052] = 249;
// bram[14053] = 252;
// bram[14054] = 253;
// bram[14055] = 253;
// bram[14056] = 251;
// bram[14057] = 248;
// bram[14058] = 243;
// bram[14059] = 236;
// bram[14060] = 228;
// bram[14061] = 219;
// bram[14062] = 208;
// bram[14063] = 196;
// bram[14064] = 183;
// bram[14065] = 170;
// bram[14066] = 156;
// bram[14067] = 142;
// bram[14068] = 127;
// bram[14069] = 112;
// bram[14070] = 98;
// bram[14071] = 84;
// bram[14072] = 70;
// bram[14073] = 58;
// bram[14074] = 46;
// bram[14075] = 35;
// bram[14076] = 25;
// bram[14077] = 17;
// bram[14078] = 11;
// bram[14079] = 5;
// bram[14080] = 2;
// bram[14081] = 0;
// bram[14082] = 0;
// bram[14083] = 1;
// bram[14084] = 4;
// bram[14085] = 9;
// bram[14086] = 15;
// bram[14087] = 23;
// bram[14088] = 32;
// bram[14089] = 43;
// bram[14090] = 54;
// bram[14091] = 67;
// bram[14092] = 80;
// bram[14093] = 94;
// bram[14094] = 108;
// bram[14095] = 123;
// bram[14096] = 138;
// bram[14097] = 152;
// bram[14098] = 166;
// bram[14099] = 180;
// bram[14100] = 193;
// bram[14101] = 205;
// bram[14102] = 216;
// bram[14103] = 226;
// bram[14104] = 234;
// bram[14105] = 241;
// bram[14106] = 247;
// bram[14107] = 251;
// bram[14108] = 253;
// bram[14109] = 253;
// bram[14110] = 252;
// bram[14111] = 250;
// bram[14112] = 245;
// bram[14113] = 239;
// bram[14114] = 232;
// bram[14115] = 223;
// bram[14116] = 213;
// bram[14117] = 201;
// bram[14118] = 189;
// bram[14119] = 176;
// bram[14120] = 162;
// bram[14121] = 148;
// bram[14122] = 133;
// bram[14123] = 118;
// bram[14124] = 104;
// bram[14125] = 90;
// bram[14126] = 76;
// bram[14127] = 63;
// bram[14128] = 51;
// bram[14129] = 39;
// bram[14130] = 29;
// bram[14131] = 21;
// bram[14132] = 13;
// bram[14133] = 7;
// bram[14134] = 3;
// bram[14135] = 0;
// bram[14136] = 0;
// bram[14137] = 0;
// bram[14138] = 3;
// bram[14139] = 7;
// bram[14140] = 12;
// bram[14141] = 20;
// bram[14142] = 28;
// bram[14143] = 38;
// bram[14144] = 49;
// bram[14145] = 61;
// bram[14146] = 74;
// bram[14147] = 88;
// bram[14148] = 102;
// bram[14149] = 117;
// bram[14150] = 131;
// bram[14151] = 146;
// bram[14152] = 160;
// bram[14153] = 174;
// bram[14154] = 188;
// bram[14155] = 200;
// bram[14156] = 211;
// bram[14157] = 222;
// bram[14158] = 231;
// bram[14159] = 238;
// bram[14160] = 245;
// bram[14161] = 249;
// bram[14162] = 252;
// bram[14163] = 253;
// bram[14164] = 253;
// bram[14165] = 251;
// bram[14166] = 247;
// bram[14167] = 242;
// bram[14168] = 235;
// bram[14169] = 227;
// bram[14170] = 217;
// bram[14171] = 206;
// bram[14172] = 194;
// bram[14173] = 181;
// bram[14174] = 168;
// bram[14175] = 154;
// bram[14176] = 139;
// bram[14177] = 125;
// bram[14178] = 110;
// bram[14179] = 96;
// bram[14180] = 82;
// bram[14181] = 68;
// bram[14182] = 56;
// bram[14183] = 44;
// bram[14184] = 33;
// bram[14185] = 24;
// bram[14186] = 16;
// bram[14187] = 10;
// bram[14188] = 5;
// bram[14189] = 1;
// bram[14190] = 0;
// bram[14191] = 0;
// bram[14192] = 1;
// bram[14193] = 5;
// bram[14194] = 10;
// bram[14195] = 16;
// bram[14196] = 24;
// bram[14197] = 34;
// bram[14198] = 44;
// bram[14199] = 56;
// bram[14200] = 69;
// bram[14201] = 82;
// bram[14202] = 96;
// bram[14203] = 111;
// bram[14204] = 125;
// bram[14205] = 140;
// bram[14206] = 154;
// bram[14207] = 168;
// bram[14208] = 182;
// bram[14209] = 195;
// bram[14210] = 207;
// bram[14211] = 217;
// bram[14212] = 227;
// bram[14213] = 235;
// bram[14214] = 242;
// bram[14215] = 247;
// bram[14216] = 251;
// bram[14217] = 253;
// bram[14218] = 253;
// bram[14219] = 252;
// bram[14220] = 249;
// bram[14221] = 244;
// bram[14222] = 238;
// bram[14223] = 230;
// bram[14224] = 221;
// bram[14225] = 211;
// bram[14226] = 199;
// bram[14227] = 187;
// bram[14228] = 174;
// bram[14229] = 160;
// bram[14230] = 145;
// bram[14231] = 131;
// bram[14232] = 116;
// bram[14233] = 102;
// bram[14234] = 87;
// bram[14235] = 74;
// bram[14236] = 61;
// bram[14237] = 49;
// bram[14238] = 38;
// bram[14239] = 28;
// bram[14240] = 19;
// bram[14241] = 12;
// bram[14242] = 7;
// bram[14243] = 3;
// bram[14244] = 0;
// bram[14245] = 0;
// bram[14246] = 1;
// bram[14247] = 3;
// bram[14248] = 8;
// bram[14249] = 13;
// bram[14250] = 21;
// bram[14251] = 30;
// bram[14252] = 40;
// bram[14253] = 51;
// bram[14254] = 63;
// bram[14255] = 77;
// bram[14256] = 90;
// bram[14257] = 105;
// bram[14258] = 119;
// bram[14259] = 134;
// bram[14260] = 148;
// bram[14261] = 163;
// bram[14262] = 176;
// bram[14263] = 190;
// bram[14264] = 202;
// bram[14265] = 213;
// bram[14266] = 223;
// bram[14267] = 232;
// bram[14268] = 239;
// bram[14269] = 245;
// bram[14270] = 250;
// bram[14271] = 252;
// bram[14272] = 253;
// bram[14273] = 253;
// bram[14274] = 250;
// bram[14275] = 246;
// bram[14276] = 241;
// bram[14277] = 234;
// bram[14278] = 225;
// bram[14279] = 215;
// bram[14280] = 204;
// bram[14281] = 192;
// bram[14282] = 179;
// bram[14283] = 166;
// bram[14284] = 151;
// bram[14285] = 137;
// bram[14286] = 122;
// bram[14287] = 108;
// bram[14288] = 93;
// bram[14289] = 79;
// bram[14290] = 66;
// bram[14291] = 54;
// bram[14292] = 42;
// bram[14293] = 32;
// bram[14294] = 23;
// bram[14295] = 15;
// bram[14296] = 9;
// bram[14297] = 4;
// bram[14298] = 1;
// bram[14299] = 0;
// bram[14300] = 0;
// bram[14301] = 2;
// bram[14302] = 6;
// bram[14303] = 11;
// bram[14304] = 18;
// bram[14305] = 26;
// bram[14306] = 35;
// bram[14307] = 46;
// bram[14308] = 58;
// bram[14309] = 71;
// bram[14310] = 84;
// bram[14311] = 99;
// bram[14312] = 113;
// bram[14313] = 128;
// bram[14314] = 142;
// bram[14315] = 157;
// bram[14316] = 171;
// bram[14317] = 184;
// bram[14318] = 197;
// bram[14319] = 208;
// bram[14320] = 219;
// bram[14321] = 228;
// bram[14322] = 237;
// bram[14323] = 243;
// bram[14324] = 248;
// bram[14325] = 252;
// bram[14326] = 253;
// bram[14327] = 253;
// bram[14328] = 252;
// bram[14329] = 248;
// bram[14330] = 243;
// bram[14331] = 237;
// bram[14332] = 229;
// bram[14333] = 220;
// bram[14334] = 209;
// bram[14335] = 197;
// bram[14336] = 185;
// bram[14337] = 171;
// bram[14338] = 158;
// bram[14339] = 143;
// bram[14340] = 128;
// bram[14341] = 114;
// bram[14342] = 99;
// bram[14343] = 85;
// bram[14344] = 72;
// bram[14345] = 59;
// bram[14346] = 47;
// bram[14347] = 36;
// bram[14348] = 26;
// bram[14349] = 18;
// bram[14350] = 11;
// bram[14351] = 6;
// bram[14352] = 2;
// bram[14353] = 0;
// bram[14354] = 0;
// bram[14355] = 1;
// bram[14356] = 4;
// bram[14357] = 8;
// bram[14358] = 15;
// bram[14359] = 22;
// bram[14360] = 31;
// bram[14361] = 42;
// bram[14362] = 53;
// bram[14363] = 65;
// bram[14364] = 79;
// bram[14365] = 93;
// bram[14366] = 107;
// bram[14367] = 121;
// bram[14368] = 136;
// bram[14369] = 151;
// bram[14370] = 165;
// bram[14371] = 178;
// bram[14372] = 191;
// bram[14373] = 204;
// bram[14374] = 215;
// bram[14375] = 225;
// bram[14376] = 233;
// bram[14377] = 241;
// bram[14378] = 246;
// bram[14379] = 250;
// bram[14380] = 253;
// bram[14381] = 253;
// bram[14382] = 253;
// bram[14383] = 250;
// bram[14384] = 246;
// bram[14385] = 240;
// bram[14386] = 233;
// bram[14387] = 224;
// bram[14388] = 214;
// bram[14389] = 203;
// bram[14390] = 190;
// bram[14391] = 177;
// bram[14392] = 163;
// bram[14393] = 149;
// bram[14394] = 135;
// bram[14395] = 120;
// bram[14396] = 105;
// bram[14397] = 91;
// bram[14398] = 77;
// bram[14399] = 64;
// bram[14400] = 52;
// bram[14401] = 41;
// bram[14402] = 30;
// bram[14403] = 21;
// bram[14404] = 14;
// bram[14405] = 8;
// bram[14406] = 3;
// bram[14407] = 1;
// bram[14408] = 0;
// bram[14409] = 0;
// bram[14410] = 2;
// bram[14411] = 6;
// bram[14412] = 12;
// bram[14413] = 19;
// bram[14414] = 27;
// bram[14415] = 37;
// bram[14416] = 48;
// bram[14417] = 60;
// bram[14418] = 73;
// bram[14419] = 87;
// bram[14420] = 101;
// bram[14421] = 115;
// bram[14422] = 130;
// bram[14423] = 144;
// bram[14424] = 159;
// bram[14425] = 173;
// bram[14426] = 186;
// bram[14427] = 199;
// bram[14428] = 210;
// bram[14429] = 221;
// bram[14430] = 230;
// bram[14431] = 238;
// bram[14432] = 244;
// bram[14433] = 249;
// bram[14434] = 252;
// bram[14435] = 253;
// bram[14436] = 253;
// bram[14437] = 251;
// bram[14438] = 248;
// bram[14439] = 243;
// bram[14440] = 236;
// bram[14441] = 228;
// bram[14442] = 218;
// bram[14443] = 207;
// bram[14444] = 196;
// bram[14445] = 183;
// bram[14446] = 169;
// bram[14447] = 155;
// bram[14448] = 141;
// bram[14449] = 126;
// bram[14450] = 112;
// bram[14451] = 97;
// bram[14452] = 83;
// bram[14453] = 70;
// bram[14454] = 57;
// bram[14455] = 45;
// bram[14456] = 34;
// bram[14457] = 25;
// bram[14458] = 17;
// bram[14459] = 10;
// bram[14460] = 5;
// bram[14461] = 2;
// bram[14462] = 0;
// bram[14463] = 0;
// bram[14464] = 1;
// bram[14465] = 4;
// bram[14466] = 9;
// bram[14467] = 16;
// bram[14468] = 24;
// bram[14469] = 33;
// bram[14470] = 43;
// bram[14471] = 55;
// bram[14472] = 67;
// bram[14473] = 81;
// bram[14474] = 95;
// bram[14475] = 109;
// bram[14476] = 124;
// bram[14477] = 138;
// bram[14478] = 153;
// bram[14479] = 167;
// bram[14480] = 181;
// bram[14481] = 193;
// bram[14482] = 205;
// bram[14483] = 216;
// bram[14484] = 226;
// bram[14485] = 235;
// bram[14486] = 241;
// bram[14487] = 247;
// bram[14488] = 251;
// bram[14489] = 253;
// bram[14490] = 253;
// bram[14491] = 252;
// bram[14492] = 249;
// bram[14493] = 245;
// bram[14494] = 239;
// bram[14495] = 231;
// bram[14496] = 222;
// bram[14497] = 212;
// bram[14498] = 201;
// bram[14499] = 188;
// bram[14500] = 175;
// bram[14501] = 161;
// bram[14502] = 147;
// bram[14503] = 132;
// bram[14504] = 118;
// bram[14505] = 103;
// bram[14506] = 89;
// bram[14507] = 75;
// bram[14508] = 62;
// bram[14509] = 50;
// bram[14510] = 39;
// bram[14511] = 29;
// bram[14512] = 20;
// bram[14513] = 13;
// bram[14514] = 7;
// bram[14515] = 3;
// bram[14516] = 0;
// bram[14517] = 0;
// bram[14518] = 0;
// bram[14519] = 3;
// bram[14520] = 7;
// bram[14521] = 13;
// bram[14522] = 20;
// bram[14523] = 29;
// bram[14524] = 39;
// bram[14525] = 50;
// bram[14526] = 62;
// bram[14527] = 75;
// bram[14528] = 89;
// bram[14529] = 103;
// bram[14530] = 118;
// bram[14531] = 132;
// bram[14532] = 147;
// bram[14533] = 161;
// bram[14534] = 175;
// bram[14535] = 188;
// bram[14536] = 201;
// bram[14537] = 212;
// bram[14538] = 222;
// bram[14539] = 231;
// bram[14540] = 239;
// bram[14541] = 245;
// bram[14542] = 249;
// bram[14543] = 252;
// bram[14544] = 253;
// bram[14545] = 253;
// bram[14546] = 251;
// bram[14547] = 247;
// bram[14548] = 242;
// bram[14549] = 235;
// bram[14550] = 226;
// bram[14551] = 217;
// bram[14552] = 206;
// bram[14553] = 194;
// bram[14554] = 181;
// bram[14555] = 167;
// bram[14556] = 153;
// bram[14557] = 139;
// bram[14558] = 124;
// bram[14559] = 109;
// bram[14560] = 95;
// bram[14561] = 81;
// bram[14562] = 68;
// bram[14563] = 55;
// bram[14564] = 43;
// bram[14565] = 33;
// bram[14566] = 24;
// bram[14567] = 16;
// bram[14568] = 9;
// bram[14569] = 4;
// bram[14570] = 1;
// bram[14571] = 0;
// bram[14572] = 0;
// bram[14573] = 2;
// bram[14574] = 5;
// bram[14575] = 10;
// bram[14576] = 17;
// bram[14577] = 25;
// bram[14578] = 34;
// bram[14579] = 45;
// bram[14580] = 57;
// bram[14581] = 69;
// bram[14582] = 83;
// bram[14583] = 97;
// bram[14584] = 111;
// bram[14585] = 126;
// bram[14586] = 141;
// bram[14587] = 155;
// bram[14588] = 169;
// bram[14589] = 183;
// bram[14590] = 195;
// bram[14591] = 207;
// bram[14592] = 218;
// bram[14593] = 228;
// bram[14594] = 236;
// bram[14595] = 242;
// bram[14596] = 248;
// bram[14597] = 251;
// bram[14598] = 253;
// bram[14599] = 253;
// bram[14600] = 252;
// bram[14601] = 249;
// bram[14602] = 244;
// bram[14603] = 238;
// bram[14604] = 230;
// bram[14605] = 221;
// bram[14606] = 210;
// bram[14607] = 199;
// bram[14608] = 186;
// bram[14609] = 173;
// bram[14610] = 159;
// bram[14611] = 145;
// bram[14612] = 130;
// bram[14613] = 115;
// bram[14614] = 101;
// bram[14615] = 87;
// bram[14616] = 73;
// bram[14617] = 60;
// bram[14618] = 48;
// bram[14619] = 37;
// bram[14620] = 27;
// bram[14621] = 19;
// bram[14622] = 12;
// bram[14623] = 6;
// bram[14624] = 2;
// bram[14625] = 0;
// bram[14626] = 0;
// bram[14627] = 1;
// bram[14628] = 3;
// bram[14629] = 8;
// bram[14630] = 14;
// bram[14631] = 21;
// bram[14632] = 30;
// bram[14633] = 40;
// bram[14634] = 52;
// bram[14635] = 64;
// bram[14636] = 77;
// bram[14637] = 91;
// bram[14638] = 105;
// bram[14639] = 120;
// bram[14640] = 134;
// bram[14641] = 149;
// bram[14642] = 163;
// bram[14643] = 177;
// bram[14644] = 190;
// bram[14645] = 202;
// bram[14646] = 214;
// bram[14647] = 224;
// bram[14648] = 232;
// bram[14649] = 240;
// bram[14650] = 246;
// bram[14651] = 250;
// bram[14652] = 253;
// bram[14653] = 253;
// bram[14654] = 253;
// bram[14655] = 250;
// bram[14656] = 246;
// bram[14657] = 241;
// bram[14658] = 233;
// bram[14659] = 225;
// bram[14660] = 215;
// bram[14661] = 204;
// bram[14662] = 192;
// bram[14663] = 179;
// bram[14664] = 165;
// bram[14665] = 151;
// bram[14666] = 136;
// bram[14667] = 122;
// bram[14668] = 107;
// bram[14669] = 93;
// bram[14670] = 79;
// bram[14671] = 66;
// bram[14672] = 53;
// bram[14673] = 42;
// bram[14674] = 31;
// bram[14675] = 22;
// bram[14676] = 15;
// bram[14677] = 8;
// bram[14678] = 4;
// bram[14679] = 1;
// bram[14680] = 0;
// bram[14681] = 0;
// bram[14682] = 2;
// bram[14683] = 6;
// bram[14684] = 11;
// bram[14685] = 18;
// bram[14686] = 26;
// bram[14687] = 36;
// bram[14688] = 47;
// bram[14689] = 59;
// bram[14690] = 72;
// bram[14691] = 85;
// bram[14692] = 99;
// bram[14693] = 114;
// bram[14694] = 128;
// bram[14695] = 143;
// bram[14696] = 157;
// bram[14697] = 171;
// bram[14698] = 185;
// bram[14699] = 197;
// bram[14700] = 209;
// bram[14701] = 220;
// bram[14702] = 229;
// bram[14703] = 237;
// bram[14704] = 243;
// bram[14705] = 248;
// bram[14706] = 252;
// bram[14707] = 253;
// bram[14708] = 253;
// bram[14709] = 252;
// bram[14710] = 248;
// bram[14711] = 243;
// bram[14712] = 237;
// bram[14713] = 229;
// bram[14714] = 219;
// bram[14715] = 209;
// bram[14716] = 197;
// bram[14717] = 184;
// bram[14718] = 171;
// bram[14719] = 157;
// bram[14720] = 142;
// bram[14721] = 128;
// bram[14722] = 113;
// bram[14723] = 99;
// bram[14724] = 85;
// bram[14725] = 71;
// bram[14726] = 58;
// bram[14727] = 46;
// bram[14728] = 36;
// bram[14729] = 26;
// bram[14730] = 18;
// bram[14731] = 11;
// bram[14732] = 6;
// bram[14733] = 2;
// bram[14734] = 0;
// bram[14735] = 0;
// bram[14736] = 1;
// bram[14737] = 4;
// bram[14738] = 9;
// bram[14739] = 15;
// bram[14740] = 23;
// bram[14741] = 32;
// bram[14742] = 42;
// bram[14743] = 54;
// bram[14744] = 66;
// bram[14745] = 79;
// bram[14746] = 93;
// bram[14747] = 108;
// bram[14748] = 122;
// bram[14749] = 137;
// bram[14750] = 151;
// bram[14751] = 165;
// bram[14752] = 179;
// bram[14753] = 192;
// bram[14754] = 204;
// bram[14755] = 215;
// bram[14756] = 225;
// bram[14757] = 234;
// bram[14758] = 241;
// bram[14759] = 246;
// bram[14760] = 250;
// bram[14761] = 253;
// bram[14762] = 253;
// bram[14763] = 252;
// bram[14764] = 250;
// bram[14765] = 245;
// bram[14766] = 240;
// bram[14767] = 232;
// bram[14768] = 223;
// bram[14769] = 213;
// bram[14770] = 202;
// bram[14771] = 190;
// bram[14772] = 177;
// bram[14773] = 163;
// bram[14774] = 149;
// bram[14775] = 134;
// bram[14776] = 119;
// bram[14777] = 105;
// bram[14778] = 90;
// bram[14779] = 77;
// bram[14780] = 64;
// bram[14781] = 51;
// bram[14782] = 40;
// bram[14783] = 30;
// bram[14784] = 21;
// bram[14785] = 14;
// bram[14786] = 8;
// bram[14787] = 3;
// bram[14788] = 1;
// bram[14789] = 0;
// bram[14790] = 0;
// bram[14791] = 2;
// bram[14792] = 6;
// bram[14793] = 12;
// bram[14794] = 19;
// bram[14795] = 28;
// bram[14796] = 38;
// bram[14797] = 49;
// bram[14798] = 61;
// bram[14799] = 74;
// bram[14800] = 87;
// bram[14801] = 101;
// bram[14802] = 116;
// bram[14803] = 131;
// bram[14804] = 145;
// bram[14805] = 160;
// bram[14806] = 173;
// bram[14807] = 187;
// bram[14808] = 199;
// bram[14809] = 211;
// bram[14810] = 221;
// bram[14811] = 230;
// bram[14812] = 238;
// bram[14813] = 244;
// bram[14814] = 249;
// bram[14815] = 252;
// bram[14816] = 253;
// bram[14817] = 253;
// bram[14818] = 251;
// bram[14819] = 247;
// bram[14820] = 242;
// bram[14821] = 235;
// bram[14822] = 227;
// bram[14823] = 218;
// bram[14824] = 207;
// bram[14825] = 195;
// bram[14826] = 182;
// bram[14827] = 169;
// bram[14828] = 155;
// bram[14829] = 140;
// bram[14830] = 126;
// bram[14831] = 111;
// bram[14832] = 96;
// bram[14833] = 82;
// bram[14834] = 69;
// bram[14835] = 56;
// bram[14836] = 45;
// bram[14837] = 34;
// bram[14838] = 25;
// bram[14839] = 17;
// bram[14840] = 10;
// bram[14841] = 5;
// bram[14842] = 1;
// bram[14843] = 0;
// bram[14844] = 0;
// bram[14845] = 1;
// bram[14846] = 5;
// bram[14847] = 10;
// bram[14848] = 16;
// bram[14849] = 24;
// bram[14850] = 33;
// bram[14851] = 44;
// bram[14852] = 55;
// bram[14853] = 68;
// bram[14854] = 81;
// bram[14855] = 95;
// bram[14856] = 110;
// bram[14857] = 124;
// bram[14858] = 139;
// bram[14859] = 154;
// bram[14860] = 168;
// bram[14861] = 181;
// bram[14862] = 194;
// bram[14863] = 206;
// bram[14864] = 217;
// bram[14865] = 227;
// bram[14866] = 235;
// bram[14867] = 242;
// bram[14868] = 247;
// bram[14869] = 251;
// bram[14870] = 253;
// bram[14871] = 253;
// bram[14872] = 252;
// bram[14873] = 249;
// bram[14874] = 245;
// bram[14875] = 239;
// bram[14876] = 231;
// bram[14877] = 222;
// bram[14878] = 212;
// bram[14879] = 200;
// bram[14880] = 188;
// bram[14881] = 174;
// bram[14882] = 161;
// bram[14883] = 146;
// bram[14884] = 132;
// bram[14885] = 117;
// bram[14886] = 103;
// bram[14887] = 88;
// bram[14888] = 75;
// bram[14889] = 62;
// bram[14890] = 49;
// bram[14891] = 38;
// bram[14892] = 28;
// bram[14893] = 20;
// bram[14894] = 13;
// bram[14895] = 7;
// bram[14896] = 3;
// bram[14897] = 0;
// bram[14898] = 0;
// bram[14899] = 0;
// bram[14900] = 3;
// bram[14901] = 7;
// bram[14902] = 13;
// bram[14903] = 20;
// bram[14904] = 29;
// bram[14905] = 39;
// bram[14906] = 50;
// bram[14907] = 63;
// bram[14908] = 76;
// bram[14909] = 89;
// bram[14910] = 104;
// bram[14911] = 118;
// bram[14912] = 133;
// bram[14913] = 147;
// bram[14914] = 162;
// bram[14915] = 176;
// bram[14916] = 189;
// bram[14917] = 201;
// bram[14918] = 212;
// bram[14919] = 223;
// bram[14920] = 232;
// bram[14921] = 239;
// bram[14922] = 245;
// bram[14923] = 250;
// bram[14924] = 252;
// bram[14925] = 253;
// bram[14926] = 253;
// bram[14927] = 251;
// bram[14928] = 247;
// bram[14929] = 241;
// bram[14930] = 234;
// bram[14931] = 226;
// bram[14932] = 216;
// bram[14933] = 205;
// bram[14934] = 193;
// bram[14935] = 180;
// bram[14936] = 167;
// bram[14937] = 152;
// bram[14938] = 138;
// bram[14939] = 123;
// bram[14940] = 109;
// bram[14941] = 94;
// bram[14942] = 80;
// bram[14943] = 67;
// bram[14944] = 54;
// bram[14945] = 43;
// bram[14946] = 32;
// bram[14947] = 23;
// bram[14948] = 15;
// bram[14949] = 9;
// bram[14950] = 4;
// bram[14951] = 1;
// bram[14952] = 0;
// bram[14953] = 0;
// bram[14954] = 2;
// bram[14955] = 5;
// bram[14956] = 10;
// bram[14957] = 17;
// bram[14958] = 25;
// bram[14959] = 35;
// bram[14960] = 46;
// bram[14961] = 57;
// bram[14962] = 70;
// bram[14963] = 84;
// bram[14964] = 98;
// bram[14965] = 112;
// bram[14966] = 127;
// bram[14967] = 141;
// bram[14968] = 156;
// bram[14969] = 170;
// bram[14970] = 183;
// bram[14971] = 196;
// bram[14972] = 208;
// bram[14973] = 218;
// bram[14974] = 228;
// bram[14975] = 236;
// bram[14976] = 243;
// bram[14977] = 248;
// bram[14978] = 251;
// bram[14979] = 253;
// bram[14980] = 253;
// bram[14981] = 252;
// bram[14982] = 249;
// bram[14983] = 244;
// bram[14984] = 237;
// bram[14985] = 230;
// bram[14986] = 220;
// bram[14987] = 210;
// bram[14988] = 198;
// bram[14989] = 186;
// bram[14990] = 172;
// bram[14991] = 158;
// bram[14992] = 144;
// bram[14993] = 129;
// bram[14994] = 115;
// bram[14995] = 100;
// bram[14996] = 86;
// bram[14997] = 73;
// bram[14998] = 60;
// bram[14999] = 48;
// bram[15000] = 37;
// bram[15001] = 27;
// bram[15002] = 19;
// bram[15003] = 12;
// bram[15004] = 6;
// bram[15005] = 2;
// bram[15006] = 0;
// bram[15007] = 0;
// bram[15008] = 1;
// bram[15009] = 4;
// bram[15010] = 8;
// bram[15011] = 14;
// bram[15012] = 22;
// bram[15013] = 31;
// bram[15014] = 41;
// bram[15015] = 52;
// bram[15016] = 65;
// bram[15017] = 78;
// bram[15018] = 92;
// bram[15019] = 106;
// bram[15020] = 121;
// bram[15021] = 135;
// bram[15022] = 150;
// bram[15023] = 164;
// bram[15024] = 178;
// bram[15025] = 191;
// bram[15026] = 203;
// bram[15027] = 214;
// bram[15028] = 224;
// bram[15029] = 233;
// bram[15030] = 240;
// bram[15031] = 246;
// bram[15032] = 250;
// bram[15033] = 253;
// bram[15034] = 253;
// bram[15035] = 253;
// bram[15036] = 250;
// bram[15037] = 246;
// bram[15038] = 240;
// bram[15039] = 233;
// bram[15040] = 224;
// bram[15041] = 214;
// bram[15042] = 203;
// bram[15043] = 191;
// bram[15044] = 178;
// bram[15045] = 164;
// bram[15046] = 150;
// bram[15047] = 136;
// bram[15048] = 121;
// bram[15049] = 106;
// bram[15050] = 92;
// bram[15051] = 78;
// bram[15052] = 65;
// bram[15053] = 53;
// bram[15054] = 41;
// bram[15055] = 31;
// bram[15056] = 22;
// bram[15057] = 14;
// bram[15058] = 8;
// bram[15059] = 4;
// bram[15060] = 1;
// bram[15061] = 0;
// bram[15062] = 0;
// bram[15063] = 2;
// bram[15064] = 6;
// bram[15065] = 11;
// bram[15066] = 18;
// bram[15067] = 27;
// bram[15068] = 36;
// bram[15069] = 47;
// bram[15070] = 59;
// bram[15071] = 72;
// bram[15072] = 86;
// bram[15073] = 100;
// bram[15074] = 114;
// bram[15075] = 129;
// bram[15076] = 144;
// bram[15077] = 158;
// bram[15078] = 172;
// bram[15079] = 185;
// bram[15080] = 198;
// bram[15081] = 210;
// bram[15082] = 220;
// bram[15083] = 229;
// bram[15084] = 237;
// bram[15085] = 244;
// bram[15086] = 249;
// bram[15087] = 252;
// bram[15088] = 253;
// bram[15089] = 253;
// bram[15090] = 251;
// bram[15091] = 248;
// bram[15092] = 243;
// bram[15093] = 236;
// bram[15094] = 228;
// bram[15095] = 219;
// bram[15096] = 208;
// bram[15097] = 196;
// bram[15098] = 184;
// bram[15099] = 170;
// bram[15100] = 156;
// bram[15101] = 142;
// bram[15102] = 127;
// bram[15103] = 112;
// bram[15104] = 98;
// bram[15105] = 84;
// bram[15106] = 70;
// bram[15107] = 58;
// bram[15108] = 46;
// bram[15109] = 35;
// bram[15110] = 26;
// bram[15111] = 17;
// bram[15112] = 11;
// bram[15113] = 5;
// bram[15114] = 2;
// bram[15115] = 0;
// bram[15116] = 0;
// bram[15117] = 1;
// bram[15118] = 4;
// bram[15119] = 9;
// bram[15120] = 15;
// bram[15121] = 23;
// bram[15122] = 32;
// bram[15123] = 43;
// bram[15124] = 54;
// bram[15125] = 67;
// bram[15126] = 80;
// bram[15127] = 94;
// bram[15128] = 108;
// bram[15129] = 123;
// bram[15130] = 137;
// bram[15131] = 152;
// bram[15132] = 166;
// bram[15133] = 180;
// bram[15134] = 193;
// bram[15135] = 205;
// bram[15136] = 216;
// bram[15137] = 226;
// bram[15138] = 234;
// bram[15139] = 241;
// bram[15140] = 247;
// bram[15141] = 251;
// bram[15142] = 253;
// bram[15143] = 253;
// bram[15144] = 252;
// bram[15145] = 250;
// bram[15146] = 245;
// bram[15147] = 239;
// bram[15148] = 232;
// bram[15149] = 223;
// bram[15150] = 213;
// bram[15151] = 201;
// bram[15152] = 189;
// bram[15153] = 176;
// bram[15154] = 162;
// bram[15155] = 148;
// bram[15156] = 133;
// bram[15157] = 119;
// bram[15158] = 104;
// bram[15159] = 90;
// bram[15160] = 76;
// bram[15161] = 63;
// bram[15162] = 51;
// bram[15163] = 39;
// bram[15164] = 29;
// bram[15165] = 21;
// bram[15166] = 13;
// bram[15167] = 7;
// bram[15168] = 3;
// bram[15169] = 0;
// bram[15170] = 0;
// bram[15171] = 0;
// bram[15172] = 3;
// bram[15173] = 7;
// bram[15174] = 12;
// bram[15175] = 20;
// bram[15176] = 28;
// bram[15177] = 38;
// bram[15178] = 49;
// bram[15179] = 61;
// bram[15180] = 74;
// bram[15181] = 88;
// bram[15182] = 102;
// bram[15183] = 117;
// bram[15184] = 131;
// bram[15185] = 146;
// bram[15186] = 160;
// bram[15187] = 174;
// bram[15188] = 187;
// bram[15189] = 200;
// bram[15190] = 211;
// bram[15191] = 222;
// bram[15192] = 231;
// bram[15193] = 238;
// bram[15194] = 245;
// bram[15195] = 249;
// bram[15196] = 252;
// bram[15197] = 253;
// bram[15198] = 253;
// bram[15199] = 251;
// bram[15200] = 247;
// bram[15201] = 242;
// bram[15202] = 235;
// bram[15203] = 227;
// bram[15204] = 217;
// bram[15205] = 206;
// bram[15206] = 194;
// bram[15207] = 182;
// bram[15208] = 168;
// bram[15209] = 154;
// bram[15210] = 139;
// bram[15211] = 125;
// bram[15212] = 110;
// bram[15213] = 96;
// bram[15214] = 82;
// bram[15215] = 68;
// bram[15216] = 56;
// bram[15217] = 44;
// bram[15218] = 34;
// bram[15219] = 24;
// bram[15220] = 16;
// bram[15221] = 10;
// bram[15222] = 5;
// bram[15223] = 1;
// bram[15224] = 0;
// bram[15225] = 0;
// bram[15226] = 1;
// bram[15227] = 5;
// bram[15228] = 10;
// bram[15229] = 16;
// bram[15230] = 24;
// bram[15231] = 34;
// bram[15232] = 44;
// bram[15233] = 56;
// bram[15234] = 69;
// bram[15235] = 82;
// bram[15236] = 96;
// bram[15237] = 110;
// bram[15238] = 125;
// bram[15239] = 140;
// bram[15240] = 154;
// bram[15241] = 168;
// bram[15242] = 182;
// bram[15243] = 195;
// bram[15244] = 207;
// bram[15245] = 217;
// bram[15246] = 227;
// bram[15247] = 235;
// bram[15248] = 242;
// bram[15249] = 247;
// bram[15250] = 251;
// bram[15251] = 253;
// bram[15252] = 253;
// bram[15253] = 252;
// bram[15254] = 249;
// bram[15255] = 244;
// bram[15256] = 238;
// bram[15257] = 230;
// bram[15258] = 221;
// bram[15259] = 211;
// bram[15260] = 200;
// bram[15261] = 187;
// bram[15262] = 174;
// bram[15263] = 160;
// bram[15264] = 146;
// bram[15265] = 131;
// bram[15266] = 116;
// bram[15267] = 102;
// bram[15268] = 88;
// bram[15269] = 74;
// bram[15270] = 61;
// bram[15271] = 49;
// bram[15272] = 38;
// bram[15273] = 28;
// bram[15274] = 19;
// bram[15275] = 12;
// bram[15276] = 7;
// bram[15277] = 3;
// bram[15278] = 0;
// bram[15279] = 0;
// bram[15280] = 1;
// bram[15281] = 3;
// bram[15282] = 7;
// bram[15283] = 13;
// bram[15284] = 21;
// bram[15285] = 30;
// bram[15286] = 40;
// bram[15287] = 51;
// bram[15288] = 63;
// bram[15289] = 76;
// bram[15290] = 90;
// bram[15291] = 104;
// bram[15292] = 119;
// bram[15293] = 134;
// bram[15294] = 148;
// bram[15295] = 162;
// bram[15296] = 176;
// bram[15297] = 189;
// bram[15298] = 202;
// bram[15299] = 213;
// bram[15300] = 223;
// bram[15301] = 232;
// bram[15302] = 239;
// bram[15303] = 245;
// bram[15304] = 250;
// bram[15305] = 252;
// bram[15306] = 253;
// bram[15307] = 253;
// bram[15308] = 251;
// bram[15309] = 247;
// bram[15310] = 241;
// bram[15311] = 234;
// bram[15312] = 225;
// bram[15313] = 216;
// bram[15314] = 204;
// bram[15315] = 192;
// bram[15316] = 179;
// bram[15317] = 166;
// bram[15318] = 152;
// bram[15319] = 137;
// bram[15320] = 123;
// bram[15321] = 108;
// bram[15322] = 94;
// bram[15323] = 80;
// bram[15324] = 66;
// bram[15325] = 54;
// bram[15326] = 42;
// bram[15327] = 32;
// bram[15328] = 23;
// bram[15329] = 15;
// bram[15330] = 9;
// bram[15331] = 4;
// bram[15332] = 1;
// bram[15333] = 0;
// bram[15334] = 0;
// bram[15335] = 2;
// bram[15336] = 5;
// bram[15337] = 11;
// bram[15338] = 17;
// bram[15339] = 26;
// bram[15340] = 35;
// bram[15341] = 46;
// bram[15342] = 58;
// bram[15343] = 71;
// bram[15344] = 84;
// bram[15345] = 98;
// bram[15346] = 113;
// bram[15347] = 127;
// bram[15348] = 142;
// bram[15349] = 156;
// bram[15350] = 170;
// bram[15351] = 184;
// bram[15352] = 197;
// bram[15353] = 208;
// bram[15354] = 219;
// bram[15355] = 228;
// bram[15356] = 236;
// bram[15357] = 243;
// bram[15358] = 248;
// bram[15359] = 251;
// bram[15360] = 253;
// bram[15361] = 253;
// bram[15362] = 252;
// bram[15363] = 248;
// bram[15364] = 244;
// bram[15365] = 237;
// bram[15366] = 229;
// bram[15367] = 220;
// bram[15368] = 209;
// bram[15369] = 198;
// bram[15370] = 185;
// bram[15371] = 172;
// bram[15372] = 158;
// bram[15373] = 143;
// bram[15374] = 129;
// bram[15375] = 114;
// bram[15376] = 100;
// bram[15377] = 85;
// bram[15378] = 72;
// bram[15379] = 59;
// bram[15380] = 47;
// bram[15381] = 36;
// bram[15382] = 27;
// bram[15383] = 18;
// bram[15384] = 11;
// bram[15385] = 6;
// bram[15386] = 2;
// bram[15387] = 0;
// bram[15388] = 0;
// bram[15389] = 1;
// bram[15390] = 4;
// bram[15391] = 8;
// bram[15392] = 14;
// bram[15393] = 22;
// bram[15394] = 31;
// bram[15395] = 41;
// bram[15396] = 53;
// bram[15397] = 65;
// bram[15398] = 78;
// bram[15399] = 92;
// bram[15400] = 107;
// bram[15401] = 121;
// bram[15402] = 136;
// bram[15403] = 150;
// bram[15404] = 165;
// bram[15405] = 178;
// bram[15406] = 191;
// bram[15407] = 203;
// bram[15408] = 215;
// bram[15409] = 225;
// bram[15410] = 233;
// bram[15411] = 240;
// bram[15412] = 246;
// bram[15413] = 250;
// bram[15414] = 253;
// bram[15415] = 253;
// bram[15416] = 253;
// bram[15417] = 250;
// bram[15418] = 246;
// bram[15419] = 240;
// bram[15420] = 233;
// bram[15421] = 224;
// bram[15422] = 214;
// bram[15423] = 203;
// bram[15424] = 190;
// bram[15425] = 177;
// bram[15426] = 164;
// bram[15427] = 149;
// bram[15428] = 135;
// bram[15429] = 120;
// bram[15430] = 106;
// bram[15431] = 91;
// bram[15432] = 78;
// bram[15433] = 64;
// bram[15434] = 52;
// bram[15435] = 41;
// bram[15436] = 30;
// bram[15437] = 22;
// bram[15438] = 14;
// bram[15439] = 8;
// bram[15440] = 3;
// bram[15441] = 1;
// bram[15442] = 0;
// bram[15443] = 0;
// bram[15444] = 2;
// bram[15445] = 6;
// bram[15446] = 12;
// bram[15447] = 19;
// bram[15448] = 27;
// bram[15449] = 37;
// bram[15450] = 48;
// bram[15451] = 60;
// bram[15452] = 73;
// bram[15453] = 86;
// bram[15454] = 101;
// bram[15455] = 115;
// bram[15456] = 130;
// bram[15457] = 144;
// bram[15458] = 159;
// bram[15459] = 173;
// bram[15460] = 186;
// bram[15461] = 198;
// bram[15462] = 210;
// bram[15463] = 221;
// bram[15464] = 230;
// bram[15465] = 238;
// bram[15466] = 244;
// bram[15467] = 249;
// bram[15468] = 252;
// bram[15469] = 253;
// bram[15470] = 253;
// bram[15471] = 251;
// bram[15472] = 248;
// bram[15473] = 243;
// bram[15474] = 236;
// bram[15475] = 228;
// bram[15476] = 218;
// bram[15477] = 208;
// bram[15478] = 196;
// bram[15479] = 183;
// bram[15480] = 170;
// bram[15481] = 155;
// bram[15482] = 141;
// bram[15483] = 126;
// bram[15484] = 112;
// bram[15485] = 97;
// bram[15486] = 83;
// bram[15487] = 70;
// bram[15488] = 57;
// bram[15489] = 45;
// bram[15490] = 35;
// bram[15491] = 25;
// bram[15492] = 17;
// bram[15493] = 10;
// bram[15494] = 5;
// bram[15495] = 2;
// bram[15496] = 0;
// bram[15497] = 0;
// bram[15498] = 1;
// bram[15499] = 4;
// bram[15500] = 9;
// bram[15501] = 16;
// bram[15502] = 23;
// bram[15503] = 33;
// bram[15504] = 43;
// bram[15505] = 55;
// bram[15506] = 67;
// bram[15507] = 81;
// bram[15508] = 95;
// bram[15509] = 109;
// bram[15510] = 124;
// bram[15511] = 138;
// bram[15512] = 153;
// bram[15513] = 167;
// bram[15514] = 180;
// bram[15515] = 193;
// bram[15516] = 205;
// bram[15517] = 216;
// bram[15518] = 226;
// bram[15519] = 234;
// bram[15520] = 241;
// bram[15521] = 247;
// bram[15522] = 251;
// bram[15523] = 253;
// bram[15524] = 253;
// bram[15525] = 252;
// bram[15526] = 249;
// bram[15527] = 245;
// bram[15528] = 239;
// bram[15529] = 231;
// bram[15530] = 222;
// bram[15531] = 212;
// bram[15532] = 201;
// bram[15533] = 188;
// bram[15534] = 175;
// bram[15535] = 161;
// bram[15536] = 147;
// bram[15537] = 133;
// bram[15538] = 118;
// bram[15539] = 103;
// bram[15540] = 89;
// bram[15541] = 75;
// bram[15542] = 62;
// bram[15543] = 50;
// bram[15544] = 39;
// bram[15545] = 29;
// bram[15546] = 20;
// bram[15547] = 13;
// bram[15548] = 7;
// bram[15549] = 3;
// bram[15550] = 0;
// bram[15551] = 0;
// bram[15552] = 0;
// bram[15553] = 3;
// bram[15554] = 7;
// bram[15555] = 13;
// bram[15556] = 20;
// bram[15557] = 29;
// bram[15558] = 39;
// bram[15559] = 50;
// bram[15560] = 62;
// bram[15561] = 75;
// bram[15562] = 89;
// bram[15563] = 103;
// bram[15564] = 117;
// bram[15565] = 132;
// bram[15566] = 147;
// bram[15567] = 161;
// bram[15568] = 175;
// bram[15569] = 188;
// bram[15570] = 200;
// bram[15571] = 212;
// bram[15572] = 222;
// bram[15573] = 231;
// bram[15574] = 239;
// bram[15575] = 245;
// bram[15576] = 249;
// bram[15577] = 252;
// bram[15578] = 253;
// bram[15579] = 253;
// bram[15580] = 251;
// bram[15581] = 247;
// bram[15582] = 242;
// bram[15583] = 235;
// bram[15584] = 226;
// bram[15585] = 217;
// bram[15586] = 206;
// bram[15587] = 194;
// bram[15588] = 181;
// bram[15589] = 167;
// bram[15590] = 153;
// bram[15591] = 139;
// bram[15592] = 124;
// bram[15593] = 109;
// bram[15594] = 95;
// bram[15595] = 81;
// bram[15596] = 68;
// bram[15597] = 55;
// bram[15598] = 44;
// bram[15599] = 33;
// bram[15600] = 24;
// bram[15601] = 16;
// bram[15602] = 9;
// bram[15603] = 5;
// bram[15604] = 1;
// bram[15605] = 0;
// bram[15606] = 0;
// bram[15607] = 2;
// bram[15608] = 5;
// bram[15609] = 10;
// bram[15610] = 17;
// bram[15611] = 25;
// bram[15612] = 34;
// bram[15613] = 45;
// bram[15614] = 57;
// bram[15615] = 69;
// bram[15616] = 83;
// bram[15617] = 97;
// bram[15618] = 111;
// bram[15619] = 126;
// bram[15620] = 140;
// bram[15621] = 155;
// bram[15622] = 169;
// bram[15623] = 182;
// bram[15624] = 195;
// bram[15625] = 207;
// bram[15626] = 218;
// bram[15627] = 227;
// bram[15628] = 236;
// bram[15629] = 242;
// bram[15630] = 248;
// bram[15631] = 251;
// bram[15632] = 253;
// bram[15633] = 253;
// bram[15634] = 252;
// bram[15635] = 249;
// bram[15636] = 244;
// bram[15637] = 238;
// bram[15638] = 230;
// bram[15639] = 221;
// bram[15640] = 210;
// bram[15641] = 199;
// bram[15642] = 186;
// bram[15643] = 173;
// bram[15644] = 159;
// bram[15645] = 145;
// bram[15646] = 130;
// bram[15647] = 116;
// bram[15648] = 101;
// bram[15649] = 87;
// bram[15650] = 73;
// bram[15651] = 60;
// bram[15652] = 48;
// bram[15653] = 37;
// bram[15654] = 28;
// bram[15655] = 19;
// bram[15656] = 12;
// bram[15657] = 6;
// bram[15658] = 2;
// bram[15659] = 0;
// bram[15660] = 0;
// bram[15661] = 1;
// bram[15662] = 3;
// bram[15663] = 8;
// bram[15664] = 14;
// bram[15665] = 21;
// bram[15666] = 30;
// bram[15667] = 40;
// bram[15668] = 52;
// bram[15669] = 64;
// bram[15670] = 77;
// bram[15671] = 91;
// bram[15672] = 105;
// bram[15673] = 120;
// bram[15674] = 134;
// bram[15675] = 149;
// bram[15676] = 163;
// bram[15677] = 177;
// bram[15678] = 190;
// bram[15679] = 202;
// bram[15680] = 213;
// bram[15681] = 224;
// bram[15682] = 232;
// bram[15683] = 240;
// bram[15684] = 246;
// bram[15685] = 250;
// bram[15686] = 253;
// bram[15687] = 253;
// bram[15688] = 253;
// bram[15689] = 250;
// bram[15690] = 246;
// bram[15691] = 241;
// bram[15692] = 234;
// bram[15693] = 225;
// bram[15694] = 215;
// bram[15695] = 204;
// bram[15696] = 192;
// bram[15697] = 179;
// bram[15698] = 165;
// bram[15699] = 151;
// bram[15700] = 136;
// bram[15701] = 122;
// bram[15702] = 107;
// bram[15703] = 93;
// bram[15704] = 79;
// bram[15705] = 66;
// bram[15706] = 53;
// bram[15707] = 42;
// bram[15708] = 32;
// bram[15709] = 22;
// bram[15710] = 15;
// bram[15711] = 9;
// bram[15712] = 4;
// bram[15713] = 1;
// bram[15714] = 0;
// bram[15715] = 0;
// bram[15716] = 2;
// bram[15717] = 6;
// bram[15718] = 11;
// bram[15719] = 18;
// bram[15720] = 26;
// bram[15721] = 36;
// bram[15722] = 47;
// bram[15723] = 59;
// bram[15724] = 71;
// bram[15725] = 85;
// bram[15726] = 99;
// bram[15727] = 113;
// bram[15728] = 128;
// bram[15729] = 143;
// bram[15730] = 157;
// bram[15731] = 171;
// bram[15732] = 185;
// bram[15733] = 197;
// bram[15734] = 209;
// bram[15735] = 219;
// bram[15736] = 229;
// bram[15737] = 237;
// bram[15738] = 243;
// bram[15739] = 248;
// bram[15740] = 252;
// bram[15741] = 253;
// bram[15742] = 253;
// bram[15743] = 252;
// bram[15744] = 248;
// bram[15745] = 243;
// bram[15746] = 237;
// bram[15747] = 229;
// bram[15748] = 219;
// bram[15749] = 209;
// bram[15750] = 197;
// bram[15751] = 184;
// bram[15752] = 171;
// bram[15753] = 157;
// bram[15754] = 143;
// bram[15755] = 128;
// bram[15756] = 113;
// bram[15757] = 99;
// bram[15758] = 85;
// bram[15759] = 71;
// bram[15760] = 58;
// bram[15761] = 47;
// bram[15762] = 36;
// bram[15763] = 26;
// bram[15764] = 18;
// bram[15765] = 11;
// bram[15766] = 6;
// bram[15767] = 2;
// bram[15768] = 0;
// bram[15769] = 0;
// bram[15770] = 1;
// bram[15771] = 4;
// bram[15772] = 9;
// bram[15773] = 15;
// bram[15774] = 22;
// bram[15775] = 32;
// bram[15776] = 42;
// bram[15777] = 53;
// bram[15778] = 66;
// bram[15779] = 79;
// bram[15780] = 93;
// bram[15781] = 107;
// bram[15782] = 122;
// bram[15783] = 137;
// bram[15784] = 151;
// bram[15785] = 165;
// bram[15786] = 179;
// bram[15787] = 192;
// bram[15788] = 204;
// bram[15789] = 215;
// bram[15790] = 225;
// bram[15791] = 234;
// bram[15792] = 241;
// bram[15793] = 246;
// bram[15794] = 250;
// bram[15795] = 253;
// bram[15796] = 253;
// bram[15797] = 253;
// bram[15798] = 250;
// bram[15799] = 246;
// bram[15800] = 240;
// bram[15801] = 232;
// bram[15802] = 223;
// bram[15803] = 213;
// bram[15804] = 202;
// bram[15805] = 190;
// bram[15806] = 177;
// bram[15807] = 163;
// bram[15808] = 149;
// bram[15809] = 134;
// bram[15810] = 120;
// bram[15811] = 105;
// bram[15812] = 91;
// bram[15813] = 77;
// bram[15814] = 64;
// bram[15815] = 51;
// bram[15816] = 40;
// bram[15817] = 30;
// bram[15818] = 21;
// bram[15819] = 14;
// bram[15820] = 8;
// bram[15821] = 3;
// bram[15822] = 1;
// bram[15823] = 0;
// bram[15824] = 0;
// bram[15825] = 2;
// bram[15826] = 6;
// bram[15827] = 12;
// bram[15828] = 19;
// bram[15829] = 28;
// bram[15830] = 37;
// bram[15831] = 48;
// bram[15832] = 60;
// bram[15833] = 73;
// bram[15834] = 87;
// bram[15835] = 101;
// bram[15836] = 116;
// bram[15837] = 130;
// bram[15838] = 145;
// bram[15839] = 159;
// bram[15840] = 173;
// bram[15841] = 187;
// bram[15842] = 199;
// bram[15843] = 211;
// bram[15844] = 221;
// bram[15845] = 230;
// bram[15846] = 238;
// bram[15847] = 244;
// bram[15848] = 249;
// bram[15849] = 252;
// bram[15850] = 253;
// bram[15851] = 253;
// bram[15852] = 251;
// bram[15853] = 248;
// bram[15854] = 242;
// bram[15855] = 236;
// bram[15856] = 227;
// bram[15857] = 218;
// bram[15858] = 207;
// bram[15859] = 195;
// bram[15860] = 182;
// bram[15861] = 169;
// bram[15862] = 155;
// bram[15863] = 140;
// bram[15864] = 126;
// bram[15865] = 111;
// bram[15866] = 97;
// bram[15867] = 83;
// bram[15868] = 69;
// bram[15869] = 57;
// bram[15870] = 45;
// bram[15871] = 34;
// bram[15872] = 25;
// bram[15873] = 17;
// bram[15874] = 10;
// bram[15875] = 5;
// bram[15876] = 2;
// bram[15877] = 0;
// bram[15878] = 0;
// bram[15879] = 1;
// bram[15880] = 5;
// bram[15881] = 9;
// bram[15882] = 16;
// bram[15883] = 24;
// bram[15884] = 33;
// bram[15885] = 44;
// bram[15886] = 55;
// bram[15887] = 68;
// bram[15888] = 81;
// bram[15889] = 95;
// bram[15890] = 110;
// bram[15891] = 124;
// bram[15892] = 139;
// bram[15893] = 153;
// bram[15894] = 167;
// bram[15895] = 181;
// bram[15896] = 194;
// bram[15897] = 206;
// bram[15898] = 217;
// bram[15899] = 226;
// bram[15900] = 235;
// bram[15901] = 242;
// bram[15902] = 247;
// bram[15903] = 251;
// bram[15904] = 253;
// bram[15905] = 253;
// bram[15906] = 252;
// bram[15907] = 249;
// bram[15908] = 245;
// bram[15909] = 239;
// bram[15910] = 231;
// bram[15911] = 222;
// bram[15912] = 212;
// bram[15913] = 200;
// bram[15914] = 188;
// bram[15915] = 175;
// bram[15916] = 161;
// bram[15917] = 146;
// bram[15918] = 132;
// bram[15919] = 117;
// bram[15920] = 103;
// bram[15921] = 88;
// bram[15922] = 75;
// bram[15923] = 62;
// bram[15924] = 50;
// bram[15925] = 38;
// bram[15926] = 29;
// bram[15927] = 20;
// bram[15928] = 13;
// bram[15929] = 7;
// bram[15930] = 3;
// bram[15931] = 0;
// bram[15932] = 0;
// bram[15933] = 0;
// bram[15934] = 3;
// bram[15935] = 7;
// bram[15936] = 13;
// bram[15937] = 20;
// bram[15938] = 29;
// bram[15939] = 39;
// bram[15940] = 50;
// bram[15941] = 62;
// bram[15942] = 76;
// bram[15943] = 89;
// bram[15944] = 103;
// bram[15945] = 118;
// bram[15946] = 133;
// bram[15947] = 147;
// bram[15948] = 162;
// bram[15949] = 175;
// bram[15950] = 189;
// bram[15951] = 201;
// bram[15952] = 212;
// bram[15953] = 222;
// bram[15954] = 231;
// bram[15955] = 239;
// bram[15956] = 245;
// bram[15957] = 249;
// bram[15958] = 252;
// bram[15959] = 253;
// bram[15960] = 253;
// bram[15961] = 251;
// bram[15962] = 247;
// bram[15963] = 241;
// bram[15964] = 234;
// bram[15965] = 226;
// bram[15966] = 216;
// bram[15967] = 205;
// bram[15968] = 193;
// bram[15969] = 180;
// bram[15970] = 167;
// bram[15971] = 153;
// bram[15972] = 138;
// bram[15973] = 123;
// bram[15974] = 109;
// bram[15975] = 94;
// bram[15976] = 80;
// bram[15977] = 67;
// bram[15978] = 55;
// bram[15979] = 43;
// bram[15980] = 33;
// bram[15981] = 23;
// bram[15982] = 15;
// bram[15983] = 9;
// bram[15984] = 4;
// bram[15985] = 1;
// bram[15986] = 0;
// bram[15987] = 0;
// bram[15988] = 2;
// bram[15989] = 5;
// bram[15990] = 10;
// bram[15991] = 17;
// bram[15992] = 25;
// bram[15993] = 35;
// bram[15994] = 45;
// bram[15995] = 57;
// bram[15996] = 70;
// bram[15997] = 83;
// bram[15998] = 97;
// bram[15999] = 112;
// bram[16000] = 127;
// bram[16001] = 143;
// bram[16002] = 159;
// bram[16003] = 175;
// bram[16004] = 189;
// bram[16005] = 203;
// bram[16006] = 215;
// bram[16007] = 226;
// bram[16008] = 236;
// bram[16009] = 243;
// bram[16010] = 249;
// bram[16011] = 252;
// bram[16012] = 253;
// bram[16013] = 253;
// bram[16014] = 250;
// bram[16015] = 245;
// bram[16016] = 238;
// bram[16017] = 229;
// bram[16018] = 219;
// bram[16019] = 207;
// bram[16020] = 194;
// bram[16021] = 179;
// bram[16022] = 164;
// bram[16023] = 148;
// bram[16024] = 132;
// bram[16025] = 115;
// bram[16026] = 99;
// bram[16027] = 83;
// bram[16028] = 68;
// bram[16029] = 54;
// bram[16030] = 41;
// bram[16031] = 30;
// bram[16032] = 20;
// bram[16033] = 12;
// bram[16034] = 6;
// bram[16035] = 2;
// bram[16036] = 0;
// bram[16037] = 0;
// bram[16038] = 2;
// bram[16039] = 6;
// bram[16040] = 12;
// bram[16041] = 21;
// bram[16042] = 31;
// bram[16043] = 42;
// bram[16044] = 55;
// bram[16045] = 69;
// bram[16046] = 84;
// bram[16047] = 100;
// bram[16048] = 116;
// bram[16049] = 133;
// bram[16050] = 149;
// bram[16051] = 165;
// bram[16052] = 180;
// bram[16053] = 194;
// bram[16054] = 208;
// bram[16055] = 220;
// bram[16056] = 230;
// bram[16057] = 239;
// bram[16058] = 245;
// bram[16059] = 250;
// bram[16060] = 253;
// bram[16061] = 253;
// bram[16062] = 252;
// bram[16063] = 248;
// bram[16064] = 243;
// bram[16065] = 235;
// bram[16066] = 226;
// bram[16067] = 215;
// bram[16068] = 202;
// bram[16069] = 189;
// bram[16070] = 174;
// bram[16071] = 158;
// bram[16072] = 142;
// bram[16073] = 126;
// bram[16074] = 109;
// bram[16075] = 93;
// bram[16076] = 78;
// bram[16077] = 63;
// bram[16078] = 49;
// bram[16079] = 37;
// bram[16080] = 26;
// bram[16081] = 17;
// bram[16082] = 10;
// bram[16083] = 4;
// bram[16084] = 1;
// bram[16085] = 0;
// bram[16086] = 0;
// bram[16087] = 3;
// bram[16088] = 8;
// bram[16089] = 15;
// bram[16090] = 24;
// bram[16091] = 35;
// bram[16092] = 47;
// bram[16093] = 60;
// bram[16094] = 75;
// bram[16095] = 90;
// bram[16096] = 106;
// bram[16097] = 122;
// bram[16098] = 139;
// bram[16099] = 155;
// bram[16100] = 170;
// bram[16101] = 185;
// bram[16102] = 199;
// bram[16103] = 212;
// bram[16104] = 224;
// bram[16105] = 233;
// bram[16106] = 241;
// bram[16107] = 247;
// bram[16108] = 251;
// bram[16109] = 253;
// bram[16110] = 253;
// bram[16111] = 251;
// bram[16112] = 247;
// bram[16113] = 240;
// bram[16114] = 232;
// bram[16115] = 222;
// bram[16116] = 210;
// bram[16117] = 197;
// bram[16118] = 183;
// bram[16119] = 168;
// bram[16120] = 152;
// bram[16121] = 136;
// bram[16122] = 120;
// bram[16123] = 103;
// bram[16124] = 87;
// bram[16125] = 72;
// bram[16126] = 58;
// bram[16127] = 45;
// bram[16128] = 33;
// bram[16129] = 23;
// bram[16130] = 14;
// bram[16131] = 7;
// bram[16132] = 3;
// bram[16133] = 0;
// bram[16134] = 0;
// bram[16135] = 1;
// bram[16136] = 5;
// bram[16137] = 11;
// bram[16138] = 18;
// bram[16139] = 28;
// bram[16140] = 39;
// bram[16141] = 51;
// bram[16142] = 65;
// bram[16143] = 80;
// bram[16144] = 96;
// bram[16145] = 112;
// bram[16146] = 128;
// bram[16147] = 145;
// bram[16148] = 161;
// bram[16149] = 176;
// bram[16150] = 191;
// bram[16151] = 204;
// bram[16152] = 217;
// bram[16153] = 227;
// bram[16154] = 236;
// bram[16155] = 244;
// bram[16156] = 249;
// bram[16157] = 252;
// bram[16158] = 253;
// bram[16159] = 253;
// bram[16160] = 250;
// bram[16161] = 244;
// bram[16162] = 237;
// bram[16163] = 228;
// bram[16164] = 218;
// bram[16165] = 206;
// bram[16166] = 192;
// bram[16167] = 178;
// bram[16168] = 162;
// bram[16169] = 146;
// bram[16170] = 130;
// bram[16171] = 114;
// bram[16172] = 97;
// bram[16173] = 82;
// bram[16174] = 67;
// bram[16175] = 53;
// bram[16176] = 40;
// bram[16177] = 29;
// bram[16178] = 19;
// bram[16179] = 11;
// bram[16180] = 5;
// bram[16181] = 1;
// bram[16182] = 0;
// bram[16183] = 0;
// bram[16184] = 2;
// bram[16185] = 7;
// bram[16186] = 13;
// bram[16187] = 22;
// bram[16188] = 32;
// bram[16189] = 43;
// bram[16190] = 56;
// bram[16191] = 71;
// bram[16192] = 86;
// bram[16193] = 102;
// bram[16194] = 118;
// bram[16195] = 134;
// bram[16196] = 150;
// bram[16197] = 166;
// bram[16198] = 182;
// bram[16199] = 196;
// bram[16200] = 209;
// bram[16201] = 221;
// bram[16202] = 231;
// bram[16203] = 239;
// bram[16204] = 246;
// bram[16205] = 250;
// bram[16206] = 253;
// bram[16207] = 253;
// bram[16208] = 252;
// bram[16209] = 248;
// bram[16210] = 242;
// bram[16211] = 234;
// bram[16212] = 225;
// bram[16213] = 214;
// bram[16214] = 201;
// bram[16215] = 187;
// bram[16216] = 172;
// bram[16217] = 156;
// bram[16218] = 140;
// bram[16219] = 124;
// bram[16220] = 108;
// bram[16221] = 92;
// bram[16222] = 76;
// bram[16223] = 62;
// bram[16224] = 48;
// bram[16225] = 36;
// bram[16226] = 25;
// bram[16227] = 16;
// bram[16228] = 9;
// bram[16229] = 4;
// bram[16230] = 1;
// bram[16231] = 0;
// bram[16232] = 1;
// bram[16233] = 4;
// bram[16234] = 9;
// bram[16235] = 16;
// bram[16236] = 25;
// bram[16237] = 36;
// bram[16238] = 48;
// bram[16239] = 61;
// bram[16240] = 76;
// bram[16241] = 91;
// bram[16242] = 108;
// bram[16243] = 124;
// bram[16244] = 140;
// bram[16245] = 156;
// bram[16246] = 172;
// bram[16247] = 187;
// bram[16248] = 201;
// bram[16249] = 213;
// bram[16250] = 225;
// bram[16251] = 234;
// bram[16252] = 242;
// bram[16253] = 248;
// bram[16254] = 252;
// bram[16255] = 253;
// bram[16256] = 253;
// bram[16257] = 251;
// bram[16258] = 246;
// bram[16259] = 239;
// bram[16260] = 231;
// bram[16261] = 221;
// bram[16262] = 209;
// bram[16263] = 196;
// bram[16264] = 182;
// bram[16265] = 166;
// bram[16266] = 151;
// bram[16267] = 134;
// bram[16268] = 118;
// bram[16269] = 102;
// bram[16270] = 86;
// bram[16271] = 71;
// bram[16272] = 56;
// bram[16273] = 43;
// bram[16274] = 32;
// bram[16275] = 22;
// bram[16276] = 13;
// bram[16277] = 7;
// bram[16278] = 2;
// bram[16279] = 0;
// bram[16280] = 0;
// bram[16281] = 1;
// bram[16282] = 5;
// bram[16283] = 11;
// bram[16284] = 19;
// bram[16285] = 29;
// bram[16286] = 40;
// bram[16287] = 53;
// bram[16288] = 67;
// bram[16289] = 82;
// bram[16290] = 97;
// bram[16291] = 114;
// bram[16292] = 130;
// bram[16293] = 146;
// bram[16294] = 162;
// bram[16295] = 178;
// bram[16296] = 192;
// bram[16297] = 206;
// bram[16298] = 218;
// bram[16299] = 228;
// bram[16300] = 237;
// bram[16301] = 244;
// bram[16302] = 249;
// bram[16303] = 253;
// bram[16304] = 253;
// bram[16305] = 252;
// bram[16306] = 249;
// bram[16307] = 244;
// bram[16308] = 237;
// bram[16309] = 227;
// bram[16310] = 217;
// bram[16311] = 204;
// bram[16312] = 191;
// bram[16313] = 176;
// bram[16314] = 161;
// bram[16315] = 145;
// bram[16316] = 128;
// bram[16317] = 112;
// bram[16318] = 96;
// bram[16319] = 80;
// bram[16320] = 65;
// bram[16321] = 51;
// bram[16322] = 39;
// bram[16323] = 28;
// bram[16324] = 18;
// bram[16325] = 11;
// bram[16326] = 5;
// bram[16327] = 1;
// bram[16328] = 0;
// bram[16329] = 0;
// bram[16330] = 3;
// bram[16331] = 7;
// bram[16332] = 14;
// bram[16333] = 23;
// bram[16334] = 33;
// bram[16335] = 45;
// bram[16336] = 58;
// bram[16337] = 72;
// bram[16338] = 87;
// bram[16339] = 103;
// bram[16340] = 120;
// bram[16341] = 136;
// bram[16342] = 152;
// bram[16343] = 168;
// bram[16344] = 183;
// bram[16345] = 197;
// bram[16346] = 210;
// bram[16347] = 222;
// bram[16348] = 232;
// bram[16349] = 240;
// bram[16350] = 246;
// bram[16351] = 251;
// bram[16352] = 253;
// bram[16353] = 253;
// bram[16354] = 251;
// bram[16355] = 247;
// bram[16356] = 241;
// bram[16357] = 233;
// bram[16358] = 224;
// bram[16359] = 212;
// bram[16360] = 200;
// bram[16361] = 186;
// bram[16362] = 171;
// bram[16363] = 155;
// bram[16364] = 139;
// bram[16365] = 122;
// bram[16366] = 106;
// bram[16367] = 90;
// bram[16368] = 75;
// bram[16369] = 60;
// bram[16370] = 47;
// bram[16371] = 35;
// bram[16372] = 24;
// bram[16373] = 15;
// bram[16374] = 8;
// bram[16375] = 3;
// bram[16376] = 0;
// bram[16377] = 0;
// bram[16378] = 1;
// bram[16379] = 4;
// bram[16380] = 10;
// bram[16381] = 17;
// bram[16382] = 26;
// bram[16383] = 37;
// bram[16384] = 49;
// bram[16385] = 63;
// bram[16386] = 78;
// bram[16387] = 93;
// bram[16388] = 109;
// bram[16389] = 126;
// bram[16390] = 142;
// bram[16391] = 158;
// bram[16392] = 174;
// bram[16393] = 188;
// bram[16394] = 202;
// bram[16395] = 215;
// bram[16396] = 226;
// bram[16397] = 235;
// bram[16398] = 243;
// bram[16399] = 248;
// bram[16400] = 252;
// bram[16401] = 253;
// bram[16402] = 253;
// bram[16403] = 250;
// bram[16404] = 245;
// bram[16405] = 239;
// bram[16406] = 230;
// bram[16407] = 220;
// bram[16408] = 208;
// bram[16409] = 195;
// bram[16410] = 180;
// bram[16411] = 165;
// bram[16412] = 149;
// bram[16413] = 133;
// bram[16414] = 116;
// bram[16415] = 100;
// bram[16416] = 84;
// bram[16417] = 69;
// bram[16418] = 55;
// bram[16419] = 42;
// bram[16420] = 31;
// bram[16421] = 21;
// bram[16422] = 12;
// bram[16423] = 6;
// bram[16424] = 2;
// bram[16425] = 0;
// bram[16426] = 0;
// bram[16427] = 2;
// bram[16428] = 6;
// bram[16429] = 12;
// bram[16430] = 20;
// bram[16431] = 30;
// bram[16432] = 41;
// bram[16433] = 54;
// bram[16434] = 68;
// bram[16435] = 83;
// bram[16436] = 99;
// bram[16437] = 115;
// bram[16438] = 132;
// bram[16439] = 148;
// bram[16440] = 164;
// bram[16441] = 179;
// bram[16442] = 194;
// bram[16443] = 207;
// bram[16444] = 219;
// bram[16445] = 229;
// bram[16446] = 238;
// bram[16447] = 245;
// bram[16448] = 250;
// bram[16449] = 253;
// bram[16450] = 253;
// bram[16451] = 252;
// bram[16452] = 249;
// bram[16453] = 243;
// bram[16454] = 236;
// bram[16455] = 226;
// bram[16456] = 215;
// bram[16457] = 203;
// bram[16458] = 189;
// bram[16459] = 175;
// bram[16460] = 159;
// bram[16461] = 143;
// bram[16462] = 127;
// bram[16463] = 110;
// bram[16464] = 94;
// bram[16465] = 79;
// bram[16466] = 64;
// bram[16467] = 50;
// bram[16468] = 38;
// bram[16469] = 27;
// bram[16470] = 17;
// bram[16471] = 10;
// bram[16472] = 4;
// bram[16473] = 1;
// bram[16474] = 0;
// bram[16475] = 0;
// bram[16476] = 3;
// bram[16477] = 8;
// bram[16478] = 15;
// bram[16479] = 23;
// bram[16480] = 34;
// bram[16481] = 46;
// bram[16482] = 59;
// bram[16483] = 74;
// bram[16484] = 89;
// bram[16485] = 105;
// bram[16486] = 121;
// bram[16487] = 138;
// bram[16488] = 154;
// bram[16489] = 170;
// bram[16490] = 185;
// bram[16491] = 199;
// bram[16492] = 212;
// bram[16493] = 223;
// bram[16494] = 233;
// bram[16495] = 241;
// bram[16496] = 247;
// bram[16497] = 251;
// bram[16498] = 253;
// bram[16499] = 253;
// bram[16500] = 251;
// bram[16501] = 247;
// bram[16502] = 241;
// bram[16503] = 232;
// bram[16504] = 223;
// bram[16505] = 211;
// bram[16506] = 198;
// bram[16507] = 184;
// bram[16508] = 169;
// bram[16509] = 153;
// bram[16510] = 137;
// bram[16511] = 121;
// bram[16512] = 104;
// bram[16513] = 88;
// bram[16514] = 73;
// bram[16515] = 59;
// bram[16516] = 45;
// bram[16517] = 33;
// bram[16518] = 23;
// bram[16519] = 14;
// bram[16520] = 8;
// bram[16521] = 3;
// bram[16522] = 0;
// bram[16523] = 0;
// bram[16524] = 1;
// bram[16525] = 5;
// bram[16526] = 10;
// bram[16527] = 18;
// bram[16528] = 27;
// bram[16529] = 38;
// bram[16530] = 51;
// bram[16531] = 64;
// bram[16532] = 79;
// bram[16533] = 95;
// bram[16534] = 111;
// bram[16535] = 127;
// bram[16536] = 144;
// bram[16537] = 160;
// bram[16538] = 175;
// bram[16539] = 190;
// bram[16540] = 204;
// bram[16541] = 216;
// bram[16542] = 227;
// bram[16543] = 236;
// bram[16544] = 243;
// bram[16545] = 249;
// bram[16546] = 252;
// bram[16547] = 253;
// bram[16548] = 253;
// bram[16549] = 250;
// bram[16550] = 245;
// bram[16551] = 238;
// bram[16552] = 229;
// bram[16553] = 218;
// bram[16554] = 206;
// bram[16555] = 193;
// bram[16556] = 179;
// bram[16557] = 163;
// bram[16558] = 147;
// bram[16559] = 131;
// bram[16560] = 115;
// bram[16561] = 98;
// bram[16562] = 83;
// bram[16563] = 68;
// bram[16564] = 54;
// bram[16565] = 41;
// bram[16566] = 29;
// bram[16567] = 20;
// bram[16568] = 12;
// bram[16569] = 6;
// bram[16570] = 2;
// bram[16571] = 0;
// bram[16572] = 0;
// bram[16573] = 2;
// bram[16574] = 6;
// bram[16575] = 13;
// bram[16576] = 21;
// bram[16577] = 31;
// bram[16578] = 43;
// bram[16579] = 56;
// bram[16580] = 70;
// bram[16581] = 85;
// bram[16582] = 101;
// bram[16583] = 117;
// bram[16584] = 133;
// bram[16585] = 150;
// bram[16586] = 165;
// bram[16587] = 181;
// bram[16588] = 195;
// bram[16589] = 208;
// bram[16590] = 220;
// bram[16591] = 230;
// bram[16592] = 239;
// bram[16593] = 246;
// bram[16594] = 250;
// bram[16595] = 253;
// bram[16596] = 253;
// bram[16597] = 252;
// bram[16598] = 248;
// bram[16599] = 242;
// bram[16600] = 235;
// bram[16601] = 225;
// bram[16602] = 214;
// bram[16603] = 202;
// bram[16604] = 188;
// bram[16605] = 173;
// bram[16606] = 157;
// bram[16607] = 141;
// bram[16608] = 125;
// bram[16609] = 109;
// bram[16610] = 93;
// bram[16611] = 77;
// bram[16612] = 62;
// bram[16613] = 49;
// bram[16614] = 36;
// bram[16615] = 26;
// bram[16616] = 17;
// bram[16617] = 9;
// bram[16618] = 4;
// bram[16619] = 1;
// bram[16620] = 0;
// bram[16621] = 0;
// bram[16622] = 3;
// bram[16623] = 9;
// bram[16624] = 16;
// bram[16625] = 24;
// bram[16626] = 35;
// bram[16627] = 47;
// bram[16628] = 61;
// bram[16629] = 75;
// bram[16630] = 91;
// bram[16631] = 107;
// bram[16632] = 123;
// bram[16633] = 139;
// bram[16634] = 155;
// bram[16635] = 171;
// bram[16636] = 186;
// bram[16637] = 200;
// bram[16638] = 213;
// bram[16639] = 224;
// bram[16640] = 234;
// bram[16641] = 242;
// bram[16642] = 248;
// bram[16643] = 251;
// bram[16644] = 253;
// bram[16645] = 253;
// bram[16646] = 251;
// bram[16647] = 246;
// bram[16648] = 240;
// bram[16649] = 232;
// bram[16650] = 221;
// bram[16651] = 210;
// bram[16652] = 197;
// bram[16653] = 183;
// bram[16654] = 167;
// bram[16655] = 152;
// bram[16656] = 135;
// bram[16657] = 119;
// bram[16658] = 103;
// bram[16659] = 87;
// bram[16660] = 72;
// bram[16661] = 57;
// bram[16662] = 44;
// bram[16663] = 32;
// bram[16664] = 22;
// bram[16665] = 14;
// bram[16666] = 7;
// bram[16667] = 3;
// bram[16668] = 0;
// bram[16669] = 0;
// bram[16670] = 1;
// bram[16671] = 5;
// bram[16672] = 11;
// bram[16673] = 19;
// bram[16674] = 28;
// bram[16675] = 39;
// bram[16676] = 52;
// bram[16677] = 66;
// bram[16678] = 81;
// bram[16679] = 96;
// bram[16680] = 113;
// bram[16681] = 129;
// bram[16682] = 145;
// bram[16683] = 161;
// bram[16684] = 177;
// bram[16685] = 191;
// bram[16686] = 205;
// bram[16687] = 217;
// bram[16688] = 228;
// bram[16689] = 237;
// bram[16690] = 244;
// bram[16691] = 249;
// bram[16692] = 252;
// bram[16693] = 253;
// bram[16694] = 252;
// bram[16695] = 249;
// bram[16696] = 244;
// bram[16697] = 237;
// bram[16698] = 228;
// bram[16699] = 217;
// bram[16700] = 205;
// bram[16701] = 192;
// bram[16702] = 177;
// bram[16703] = 162;
// bram[16704] = 146;
// bram[16705] = 129;
// bram[16706] = 113;
// bram[16707] = 97;
// bram[16708] = 81;
// bram[16709] = 66;
// bram[16710] = 52;
// bram[16711] = 40;
// bram[16712] = 28;
// bram[16713] = 19;
// bram[16714] = 11;
// bram[16715] = 5;
// bram[16716] = 1;
// bram[16717] = 0;
// bram[16718] = 0;
// bram[16719] = 2;
// bram[16720] = 7;
// bram[16721] = 14;
// bram[16722] = 22;
// bram[16723] = 32;
// bram[16724] = 44;
// bram[16725] = 57;
// bram[16726] = 71;
// bram[16727] = 86;
// bram[16728] = 102;
// bram[16729] = 119;
// bram[16730] = 135;
// bram[16731] = 151;
// bram[16732] = 167;
// bram[16733] = 182;
// bram[16734] = 196;
// bram[16735] = 210;
// bram[16736] = 221;
// bram[16737] = 231;
// bram[16738] = 240;
// bram[16739] = 246;
// bram[16740] = 251;
// bram[16741] = 253;
// bram[16742] = 253;
// bram[16743] = 252;
// bram[16744] = 248;
// bram[16745] = 242;
// bram[16746] = 234;
// bram[16747] = 224;
// bram[16748] = 213;
// bram[16749] = 200;
// bram[16750] = 186;
// bram[16751] = 171;
// bram[16752] = 156;
// bram[16753] = 140;
// bram[16754] = 123;
// bram[16755] = 107;
// bram[16756] = 91;
// bram[16757] = 75;
// bram[16758] = 61;
// bram[16759] = 47;
// bram[16760] = 35;
// bram[16761] = 25;
// bram[16762] = 16;
// bram[16763] = 9;
// bram[16764] = 4;
// bram[16765] = 0;
// bram[16766] = 0;
// bram[16767] = 1;
// bram[16768] = 4;
// bram[16769] = 9;
// bram[16770] = 16;
// bram[16771] = 26;
// bram[16772] = 36;
// bram[16773] = 49;
// bram[16774] = 62;
// bram[16775] = 77;
// bram[16776] = 92;
// bram[16777] = 108;
// bram[16778] = 125;
// bram[16779] = 141;
// bram[16780] = 157;
// bram[16781] = 173;
// bram[16782] = 188;
// bram[16783] = 201;
// bram[16784] = 214;
// bram[16785] = 225;
// bram[16786] = 235;
// bram[16787] = 242;
// bram[16788] = 248;
// bram[16789] = 252;
// bram[16790] = 253;
// bram[16791] = 253;
// bram[16792] = 250;
// bram[16793] = 246;
// bram[16794] = 239;
// bram[16795] = 231;
// bram[16796] = 220;
// bram[16797] = 208;
// bram[16798] = 195;
// bram[16799] = 181;
// bram[16800] = 166;
// bram[16801] = 150;
// bram[16802] = 134;
// bram[16803] = 117;
// bram[16804] = 101;
// bram[16805] = 85;
// bram[16806] = 70;
// bram[16807] = 56;
// bram[16808] = 43;
// bram[16809] = 31;
// bram[16810] = 21;
// bram[16811] = 13;
// bram[16812] = 7;
// bram[16813] = 2;
// bram[16814] = 0;
// bram[16815] = 0;
// bram[16816] = 2;
// bram[16817] = 6;
// bram[16818] = 12;
// bram[16819] = 20;
// bram[16820] = 29;
// bram[16821] = 41;
// bram[16822] = 53;
// bram[16823] = 67;
// bram[16824] = 82;
// bram[16825] = 98;
// bram[16826] = 114;
// bram[16827] = 131;
// bram[16828] = 147;
// bram[16829] = 163;
// bram[16830] = 178;
// bram[16831] = 193;
// bram[16832] = 206;
// bram[16833] = 218;
// bram[16834] = 229;
// bram[16835] = 238;
// bram[16836] = 245;
// bram[16837] = 250;
// bram[16838] = 253;
// bram[16839] = 253;
// bram[16840] = 252;
// bram[16841] = 249;
// bram[16842] = 243;
// bram[16843] = 236;
// bram[16844] = 227;
// bram[16845] = 216;
// bram[16846] = 204;
// bram[16847] = 190;
// bram[16848] = 175;
// bram[16849] = 160;
// bram[16850] = 144;
// bram[16851] = 128;
// bram[16852] = 111;
// bram[16853] = 95;
// bram[16854] = 79;
// bram[16855] = 65;
// bram[16856] = 51;
// bram[16857] = 38;
// bram[16858] = 27;
// bram[16859] = 18;
// bram[16860] = 10;
// bram[16861] = 5;
// bram[16862] = 1;
// bram[16863] = 0;
// bram[16864] = 0;
// bram[16865] = 3;
// bram[16866] = 8;
// bram[16867] = 14;
// bram[16868] = 23;
// bram[16869] = 33;
// bram[16870] = 45;
// bram[16871] = 58;
// bram[16872] = 73;
// bram[16873] = 88;
// bram[16874] = 104;
// bram[16875] = 120;
// bram[16876] = 137;
// bram[16877] = 153;
// bram[16878] = 169;
// bram[16879] = 184;
// bram[16880] = 198;
// bram[16881] = 211;
// bram[16882] = 222;
// bram[16883] = 232;
// bram[16884] = 240;
// bram[16885] = 247;
// bram[16886] = 251;
// bram[16887] = 253;
// bram[16888] = 253;
// bram[16889] = 251;
// bram[16890] = 247;
// bram[16891] = 241;
// bram[16892] = 233;
// bram[16893] = 223;
// bram[16894] = 212;
// bram[16895] = 199;
// bram[16896] = 185;
// bram[16897] = 170;
// bram[16898] = 154;
// bram[16899] = 138;
// bram[16900] = 122;
// bram[16901] = 105;
// bram[16902] = 89;
// bram[16903] = 74;
// bram[16904] = 59;
// bram[16905] = 46;
// bram[16906] = 34;
// bram[16907] = 24;
// bram[16908] = 15;
// bram[16909] = 8;
// bram[16910] = 3;
// bram[16911] = 0;
// bram[16912] = 0;
// bram[16913] = 1;
// bram[16914] = 4;
// bram[16915] = 10;
// bram[16916] = 17;
// bram[16917] = 27;
// bram[16918] = 37;
// bram[16919] = 50;
// bram[16920] = 64;
// bram[16921] = 78;
// bram[16922] = 94;
// bram[16923] = 110;
// bram[16924] = 126;
// bram[16925] = 143;
// bram[16926] = 159;
// bram[16927] = 174;
// bram[16928] = 189;
// bram[16929] = 203;
// bram[16930] = 215;
// bram[16931] = 226;
// bram[16932] = 236;
// bram[16933] = 243;
// bram[16934] = 249;
// bram[16935] = 252;
// bram[16936] = 253;
// bram[16937] = 253;
// bram[16938] = 250;
// bram[16939] = 245;
// bram[16940] = 238;
// bram[16941] = 230;
// bram[16942] = 219;
// bram[16943] = 207;
// bram[16944] = 194;
// bram[16945] = 179;
// bram[16946] = 164;
// bram[16947] = 148;
// bram[16948] = 132;
// bram[16949] = 115;
// bram[16950] = 99;
// bram[16951] = 84;
// bram[16952] = 68;
// bram[16953] = 54;
// bram[16954] = 42;
// bram[16955] = 30;
// bram[16956] = 20;
// bram[16957] = 12;
// bram[16958] = 6;
// bram[16959] = 2;
// bram[16960] = 0;
// bram[16961] = 0;
// bram[16962] = 2;
// bram[16963] = 6;
// bram[16964] = 12;
// bram[16965] = 20;
// bram[16966] = 30;
// bram[16967] = 42;
// bram[16968] = 55;
// bram[16969] = 69;
// bram[16970] = 84;
// bram[16971] = 100;
// bram[16972] = 116;
// bram[16973] = 132;
// bram[16974] = 149;
// bram[16975] = 165;
// bram[16976] = 180;
// bram[16977] = 194;
// bram[16978] = 208;
// bram[16979] = 219;
// bram[16980] = 230;
// bram[16981] = 238;
// bram[16982] = 245;
// bram[16983] = 250;
// bram[16984] = 253;
// bram[16985] = 253;
// bram[16986] = 252;
// bram[16987] = 248;
// bram[16988] = 243;
// bram[16989] = 235;
// bram[16990] = 226;
// bram[16991] = 215;
// bram[16992] = 202;
// bram[16993] = 189;
// bram[16994] = 174;
// bram[16995] = 158;
// bram[16996] = 142;
// bram[16997] = 126;
// bram[16998] = 109;
// bram[16999] = 93;
// bram[17000] = 78;
// bram[17001] = 63;
// bram[17002] = 50;
// bram[17003] = 37;
// bram[17004] = 26;
// bram[17005] = 17;
// bram[17006] = 10;
// bram[17007] = 4;
// bram[17008] = 1;
// bram[17009] = 0;
// bram[17010] = 0;
// bram[17011] = 3;
// bram[17012] = 8;
// bram[17013] = 15;
// bram[17014] = 24;
// bram[17015] = 34;
// bram[17016] = 46;
// bram[17017] = 60;
// bram[17018] = 74;
// bram[17019] = 90;
// bram[17020] = 106;
// bram[17021] = 122;
// bram[17022] = 138;
// bram[17023] = 155;
// bram[17024] = 170;
// bram[17025] = 185;
// bram[17026] = 199;
// bram[17027] = 212;
// bram[17028] = 223;
// bram[17029] = 233;
// bram[17030] = 241;
// bram[17031] = 247;
// bram[17032] = 251;
// bram[17033] = 253;
// bram[17034] = 253;
// bram[17035] = 251;
// bram[17036] = 247;
// bram[17037] = 240;
// bram[17038] = 232;
// bram[17039] = 222;
// bram[17040] = 210;
// bram[17041] = 198;
// bram[17042] = 183;
// bram[17043] = 168;
// bram[17044] = 152;
// bram[17045] = 136;
// bram[17046] = 120;
// bram[17047] = 104;
// bram[17048] = 88;
// bram[17049] = 72;
// bram[17050] = 58;
// bram[17051] = 45;
// bram[17052] = 33;
// bram[17053] = 23;
// bram[17054] = 14;
// bram[17055] = 7;
// bram[17056] = 3;
// bram[17057] = 0;
// bram[17058] = 0;
// bram[17059] = 1;
// bram[17060] = 5;
// bram[17061] = 11;
// bram[17062] = 18;
// bram[17063] = 28;
// bram[17064] = 39;
// bram[17065] = 51;
// bram[17066] = 65;
// bram[17067] = 80;
// bram[17068] = 95;
// bram[17069] = 112;
// bram[17070] = 128;
// bram[17071] = 144;
// bram[17072] = 160;
// bram[17073] = 176;
// bram[17074] = 191;
// bram[17075] = 204;
// bram[17076] = 216;
// bram[17077] = 227;
// bram[17078] = 236;
// bram[17079] = 244;
// bram[17080] = 249;
// bram[17081] = 252;
// bram[17082] = 253;
// bram[17083] = 253;
// bram[17084] = 250;
// bram[17085] = 244;
// bram[17086] = 237;
// bram[17087] = 229;
// bram[17088] = 218;
// bram[17089] = 206;
// bram[17090] = 192;
// bram[17091] = 178;
// bram[17092] = 163;
// bram[17093] = 147;
// bram[17094] = 130;
// bram[17095] = 114;
// bram[17096] = 98;
// bram[17097] = 82;
// bram[17098] = 67;
// bram[17099] = 53;
// bram[17100] = 40;
// bram[17101] = 29;
// bram[17102] = 19;
// bram[17103] = 11;
// bram[17104] = 5;
// bram[17105] = 2;
// bram[17106] = 0;
// bram[17107] = 0;
// bram[17108] = 2;
// bram[17109] = 7;
// bram[17110] = 13;
// bram[17111] = 21;
// bram[17112] = 32;
// bram[17113] = 43;
// bram[17114] = 56;
// bram[17115] = 70;
// bram[17116] = 86;
// bram[17117] = 101;
// bram[17118] = 118;
// bram[17119] = 134;
// bram[17120] = 150;
// bram[17121] = 166;
// bram[17122] = 181;
// bram[17123] = 196;
// bram[17124] = 209;
// bram[17125] = 221;
// bram[17126] = 231;
// bram[17127] = 239;
// bram[17128] = 246;
// bram[17129] = 250;
// bram[17130] = 253;
// bram[17131] = 253;
// bram[17132] = 252;
// bram[17133] = 248;
// bram[17134] = 242;
// bram[17135] = 234;
// bram[17136] = 225;
// bram[17137] = 214;
// bram[17138] = 201;
// bram[17139] = 187;
// bram[17140] = 172;
// bram[17141] = 157;
// bram[17142] = 141;
// bram[17143] = 124;
// bram[17144] = 108;
// bram[17145] = 92;
// bram[17146] = 76;
// bram[17147] = 62;
// bram[17148] = 48;
// bram[17149] = 36;
// bram[17150] = 25;
// bram[17151] = 16;
// bram[17152] = 9;
// bram[17153] = 4;
// bram[17154] = 1;
// bram[17155] = 0;
// bram[17156] = 1;
// bram[17157] = 4;
// bram[17158] = 9;
// bram[17159] = 16;
// bram[17160] = 25;
// bram[17161] = 36;
// bram[17162] = 48;
// bram[17163] = 61;
// bram[17164] = 76;
// bram[17165] = 91;
// bram[17166] = 107;
// bram[17167] = 124;
// bram[17168] = 140;
// bram[17169] = 156;
// bram[17170] = 172;
// bram[17171] = 187;
// bram[17172] = 201;
// bram[17173] = 213;
// bram[17174] = 225;
// bram[17175] = 234;
// bram[17176] = 242;
// bram[17177] = 248;
// bram[17178] = 252;
// bram[17179] = 253;
// bram[17180] = 253;
// bram[17181] = 251;
// bram[17182] = 246;
// bram[17183] = 239;
// bram[17184] = 231;
// bram[17185] = 221;
// bram[17186] = 209;
// bram[17187] = 196;
// bram[17188] = 182;
// bram[17189] = 167;
// bram[17190] = 151;
// bram[17191] = 135;
// bram[17192] = 118;
// bram[17193] = 102;
// bram[17194] = 86;
// bram[17195] = 71;
// bram[17196] = 57;
// bram[17197] = 44;
// bram[17198] = 32;
// bram[17199] = 22;
// bram[17200] = 13;
// bram[17201] = 7;
// bram[17202] = 2;
// bram[17203] = 0;
// bram[17204] = 0;
// bram[17205] = 1;
// bram[17206] = 5;
// bram[17207] = 11;
// bram[17208] = 19;
// bram[17209] = 29;
// bram[17210] = 40;
// bram[17211] = 53;
// bram[17212] = 67;
// bram[17213] = 81;
// bram[17214] = 97;
// bram[17215] = 113;
// bram[17216] = 130;
// bram[17217] = 146;
// bram[17218] = 162;
// bram[17219] = 177;
// bram[17220] = 192;
// bram[17221] = 205;
// bram[17222] = 218;
// bram[17223] = 228;
// bram[17224] = 237;
// bram[17225] = 244;
// bram[17226] = 249;
// bram[17227] = 253;
// bram[17228] = 253;
// bram[17229] = 252;
// bram[17230] = 249;
// bram[17231] = 244;
// bram[17232] = 237;
// bram[17233] = 228;
// bram[17234] = 217;
// bram[17235] = 205;
// bram[17236] = 191;
// bram[17237] = 176;
// bram[17238] = 161;
// bram[17239] = 145;
// bram[17240] = 128;
// bram[17241] = 112;
// bram[17242] = 96;
// bram[17243] = 80;
// bram[17244] = 65;
// bram[17245] = 52;
// bram[17246] = 39;
// bram[17247] = 28;
// bram[17248] = 18;
// bram[17249] = 11;
// bram[17250] = 5;
// bram[17251] = 1;
// bram[17252] = 0;
// bram[17253] = 0;
// bram[17254] = 3;
// bram[17255] = 7;
// bram[17256] = 14;
// bram[17257] = 22;
// bram[17258] = 33;
// bram[17259] = 44;
// bram[17260] = 58;
// bram[17261] = 72;
// bram[17262] = 87;
// bram[17263] = 103;
// bram[17264] = 119;
// bram[17265] = 136;
// bram[17266] = 152;
// bram[17267] = 168;
// bram[17268] = 183;
// bram[17269] = 197;
// bram[17270] = 210;
// bram[17271] = 222;
// bram[17272] = 232;
// bram[17273] = 240;
// bram[17274] = 246;
// bram[17275] = 251;
// bram[17276] = 253;
// bram[17277] = 253;
// bram[17278] = 251;
// bram[17279] = 247;
// bram[17280] = 241;
// bram[17281] = 233;
// bram[17282] = 224;
// bram[17283] = 212;
// bram[17284] = 200;
// bram[17285] = 186;
// bram[17286] = 171;
// bram[17287] = 155;
// bram[17288] = 139;
// bram[17289] = 122;
// bram[17290] = 106;
// bram[17291] = 90;
// bram[17292] = 75;
// bram[17293] = 60;
// bram[17294] = 47;
// bram[17295] = 35;
// bram[17296] = 24;
// bram[17297] = 15;
// bram[17298] = 8;
// bram[17299] = 3;
// bram[17300] = 0;
// bram[17301] = 0;
// bram[17302] = 1;
// bram[17303] = 4;
// bram[17304] = 9;
// bram[17305] = 17;
// bram[17306] = 26;
// bram[17307] = 37;
// bram[17308] = 49;
// bram[17309] = 63;
// bram[17310] = 77;
// bram[17311] = 93;
// bram[17312] = 109;
// bram[17313] = 125;
// bram[17314] = 142;
// bram[17315] = 158;
// bram[17316] = 173;
// bram[17317] = 188;
// bram[17318] = 202;
// bram[17319] = 215;
// bram[17320] = 226;
// bram[17321] = 235;
// bram[17322] = 243;
// bram[17323] = 248;
// bram[17324] = 252;
// bram[17325] = 253;
// bram[17326] = 253;
// bram[17327] = 250;
// bram[17328] = 245;
// bram[17329] = 239;
// bram[17330] = 230;
// bram[17331] = 220;
// bram[17332] = 208;
// bram[17333] = 195;
// bram[17334] = 180;
// bram[17335] = 165;
// bram[17336] = 149;
// bram[17337] = 133;
// bram[17338] = 116;
// bram[17339] = 100;
// bram[17340] = 84;
// bram[17341] = 69;
// bram[17342] = 55;
// bram[17343] = 42;
// bram[17344] = 31;
// bram[17345] = 21;
// bram[17346] = 13;
// bram[17347] = 6;
// bram[17348] = 2;
// bram[17349] = 0;
// bram[17350] = 0;
// bram[17351] = 2;
// bram[17352] = 6;
// bram[17353] = 12;
// bram[17354] = 20;
// bram[17355] = 30;
// bram[17356] = 41;
// bram[17357] = 54;
// bram[17358] = 68;
// bram[17359] = 83;
// bram[17360] = 99;
// bram[17361] = 115;
// bram[17362] = 131;
// bram[17363] = 148;
// bram[17364] = 164;
// bram[17365] = 179;
// bram[17366] = 193;
// bram[17367] = 207;
// bram[17368] = 219;
// bram[17369] = 229;
// bram[17370] = 238;
// bram[17371] = 245;
// bram[17372] = 250;
// bram[17373] = 253;
// bram[17374] = 253;
// bram[17375] = 252;
// bram[17376] = 249;
// bram[17377] = 243;
// bram[17378] = 236;
// bram[17379] = 227;
// bram[17380] = 216;
// bram[17381] = 203;
// bram[17382] = 190;
// bram[17383] = 175;
// bram[17384] = 159;
// bram[17385] = 143;
// bram[17386] = 127;
// bram[17387] = 110;
// bram[17388] = 94;
// bram[17389] = 79;
// bram[17390] = 64;
// bram[17391] = 50;
// bram[17392] = 38;
// bram[17393] = 27;
// bram[17394] = 18;
// bram[17395] = 10;
// bram[17396] = 4;
// bram[17397] = 1;
// bram[17398] = 0;
// bram[17399] = 0;
// bram[17400] = 3;
// bram[17401] = 8;
// bram[17402] = 15;
// bram[17403] = 23;
// bram[17404] = 34;
// bram[17405] = 46;
// bram[17406] = 59;
// bram[17407] = 73;
// bram[17408] = 89;
// bram[17409] = 105;
// bram[17410] = 121;
// bram[17411] = 137;
// bram[17412] = 154;
// bram[17413] = 169;
// bram[17414] = 184;
// bram[17415] = 199;
// bram[17416] = 211;
// bram[17417] = 223;
// bram[17418] = 233;
// bram[17419] = 241;
// bram[17420] = 247;
// bram[17421] = 251;
// bram[17422] = 253;
// bram[17423] = 253;
// bram[17424] = 251;
// bram[17425] = 247;
// bram[17426] = 241;
// bram[17427] = 233;
// bram[17428] = 223;
// bram[17429] = 211;
// bram[17430] = 198;
// bram[17431] = 184;
// bram[17432] = 169;
// bram[17433] = 153;
// bram[17434] = 137;
// bram[17435] = 121;
// bram[17436] = 104;
// bram[17437] = 89;
// bram[17438] = 73;
// bram[17439] = 59;
// bram[17440] = 46;
// bram[17441] = 34;
// bram[17442] = 23;
// bram[17443] = 15;
// bram[17444] = 8;
// bram[17445] = 3;
// bram[17446] = 0;
// bram[17447] = 0;
// bram[17448] = 1;
// bram[17449] = 5;
// bram[17450] = 10;
// bram[17451] = 18;
// bram[17452] = 27;
// bram[17453] = 38;
// bram[17454] = 50;
// bram[17455] = 64;
// bram[17456] = 79;
// bram[17457] = 95;
// bram[17458] = 111;
// bram[17459] = 127;
// bram[17460] = 143;
// bram[17461] = 159;
// bram[17462] = 175;
// bram[17463] = 190;
// bram[17464] = 203;
// bram[17465] = 216;
// bram[17466] = 227;
// bram[17467] = 236;
// bram[17468] = 243;
// bram[17469] = 249;
// bram[17470] = 252;
// bram[17471] = 253;
// bram[17472] = 253;
// bram[17473] = 250;
// bram[17474] = 245;
// bram[17475] = 238;
// bram[17476] = 229;
// bram[17477] = 219;
// bram[17478] = 207;
// bram[17479] = 193;
// bram[17480] = 179;
// bram[17481] = 163;
// bram[17482] = 147;
// bram[17483] = 131;
// bram[17484] = 115;
// bram[17485] = 99;
// bram[17486] = 83;
// bram[17487] = 68;
// bram[17488] = 54;
// bram[17489] = 41;
// bram[17490] = 30;
// bram[17491] = 20;
// bram[17492] = 12;
// bram[17493] = 6;
// bram[17494] = 2;
// bram[17495] = 0;
// bram[17496] = 0;
// bram[17497] = 2;
// bram[17498] = 6;
// bram[17499] = 13;
// bram[17500] = 21;
// bram[17501] = 31;
// bram[17502] = 42;
// bram[17503] = 55;
// bram[17504] = 70;
// bram[17505] = 85;
// bram[17506] = 100;
// bram[17507] = 117;
// bram[17508] = 133;
// bram[17509] = 149;
// bram[17510] = 165;
// bram[17511] = 181;
// bram[17512] = 195;
// bram[17513] = 208;
// bram[17514] = 220;
// bram[17515] = 230;
// bram[17516] = 239;
// bram[17517] = 246;
// bram[17518] = 250;
// bram[17519] = 253;
// bram[17520] = 253;
// bram[17521] = 252;
// bram[17522] = 248;
// bram[17523] = 243;
// bram[17524] = 235;
// bram[17525] = 225;
// bram[17526] = 214;
// bram[17527] = 202;
// bram[17528] = 188;
// bram[17529] = 173;
// bram[17530] = 158;
// bram[17531] = 141;
// bram[17532] = 125;
// bram[17533] = 109;
// bram[17534] = 93;
// bram[17535] = 77;
// bram[17536] = 63;
// bram[17537] = 49;
// bram[17538] = 37;
// bram[17539] = 26;
// bram[17540] = 17;
// bram[17541] = 9;
// bram[17542] = 4;
// bram[17543] = 1;
// bram[17544] = 0;
// bram[17545] = 0;
// bram[17546] = 3;
// bram[17547] = 8;
// bram[17548] = 15;
// bram[17549] = 24;
// bram[17550] = 35;
// bram[17551] = 47;
// bram[17552] = 60;
// bram[17553] = 75;
// bram[17554] = 90;
// bram[17555] = 106;
// bram[17556] = 123;
// bram[17557] = 139;
// bram[17558] = 155;
// bram[17559] = 171;
// bram[17560] = 186;
// bram[17561] = 200;
// bram[17562] = 213;
// bram[17563] = 224;
// bram[17564] = 234;
// bram[17565] = 242;
// bram[17566] = 247;
// bram[17567] = 251;
// bram[17568] = 253;
// bram[17569] = 253;
// bram[17570] = 251;
// bram[17571] = 246;
// bram[17572] = 240;
// bram[17573] = 232;
// bram[17574] = 222;
// bram[17575] = 210;
// bram[17576] = 197;
// bram[17577] = 183;
// bram[17578] = 168;
// bram[17579] = 152;
// bram[17580] = 135;
// bram[17581] = 119;
// bram[17582] = 103;
// bram[17583] = 87;
// bram[17584] = 72;
// bram[17585] = 57;
// bram[17586] = 44;
// bram[17587] = 32;
// bram[17588] = 22;
// bram[17589] = 14;
// bram[17590] = 7;
// bram[17591] = 3;
// bram[17592] = 0;
// bram[17593] = 0;
// bram[17594] = 1;
// bram[17595] = 5;
// bram[17596] = 11;
// bram[17597] = 19;
// bram[17598] = 28;
// bram[17599] = 39;
// bram[17600] = 52;
// bram[17601] = 66;
// bram[17602] = 81;
// bram[17603] = 96;
// bram[17604] = 112;
// bram[17605] = 129;
// bram[17606] = 145;
// bram[17607] = 161;
// bram[17608] = 177;
// bram[17609] = 191;
// bram[17610] = 205;
// bram[17611] = 217;
// bram[17612] = 228;
// bram[17613] = 237;
// bram[17614] = 244;
// bram[17615] = 249;
// bram[17616] = 252;
// bram[17617] = 253;
// bram[17618] = 252;
// bram[17619] = 249;
// bram[17620] = 244;
// bram[17621] = 237;
// bram[17622] = 228;
// bram[17623] = 217;
// bram[17624] = 205;
// bram[17625] = 192;
// bram[17626] = 177;
// bram[17627] = 162;
// bram[17628] = 146;
// bram[17629] = 129;
// bram[17630] = 113;
// bram[17631] = 97;
// bram[17632] = 81;
// bram[17633] = 66;
// bram[17634] = 52;
// bram[17635] = 40;
// bram[17636] = 29;
// bram[17637] = 19;
// bram[17638] = 11;
// bram[17639] = 5;
// bram[17640] = 1;
// bram[17641] = 0;
// bram[17642] = 0;
// bram[17643] = 2;
// bram[17644] = 7;
// bram[17645] = 13;
// bram[17646] = 22;
// bram[17647] = 32;
// bram[17648] = 44;
// bram[17649] = 57;
// bram[17650] = 71;
// bram[17651] = 86;
// bram[17652] = 102;
// bram[17653] = 118;
// bram[17654] = 135;
// bram[17655] = 151;
// bram[17656] = 167;
// bram[17657] = 182;
// bram[17658] = 196;
// bram[17659] = 209;
// bram[17660] = 221;
// bram[17661] = 231;
// bram[17662] = 240;
// bram[17663] = 246;
// bram[17664] = 251;
// bram[17665] = 253;
// bram[17666] = 253;
// bram[17667] = 252;
// bram[17668] = 248;
// bram[17669] = 242;
// bram[17670] = 234;
// bram[17671] = 224;
// bram[17672] = 213;
// bram[17673] = 200;
// bram[17674] = 187;
// bram[17675] = 172;
// bram[17676] = 156;
// bram[17677] = 140;
// bram[17678] = 123;
// bram[17679] = 107;
// bram[17680] = 91;
// bram[17681] = 76;
// bram[17682] = 61;
// bram[17683] = 48;
// bram[17684] = 35;
// bram[17685] = 25;
// bram[17686] = 16;
// bram[17687] = 9;
// bram[17688] = 4;
// bram[17689] = 0;
// bram[17690] = 0;
// bram[17691] = 1;
// bram[17692] = 4;
// bram[17693] = 9;
// bram[17694] = 16;
// bram[17695] = 25;
// bram[17696] = 36;
// bram[17697] = 48;
// bram[17698] = 62;
// bram[17699] = 77;
// bram[17700] = 92;
// bram[17701] = 108;
// bram[17702] = 124;
// bram[17703] = 141;
// bram[17704] = 157;
// bram[17705] = 173;
// bram[17706] = 187;
// bram[17707] = 201;
// bram[17708] = 214;
// bram[17709] = 225;
// bram[17710] = 235;
// bram[17711] = 242;
// bram[17712] = 248;
// bram[17713] = 252;
// bram[17714] = 253;
// bram[17715] = 253;
// bram[17716] = 250;
// bram[17717] = 246;
// bram[17718] = 239;
// bram[17719] = 231;
// bram[17720] = 220;
// bram[17721] = 209;
// bram[17722] = 195;
// bram[17723] = 181;
// bram[17724] = 166;
// bram[17725] = 150;
// bram[17726] = 134;
// bram[17727] = 117;
// bram[17728] = 101;
// bram[17729] = 85;
// bram[17730] = 70;
// bram[17731] = 56;
// bram[17732] = 43;
// bram[17733] = 31;
// bram[17734] = 21;
// bram[17735] = 13;
// bram[17736] = 7;
// bram[17737] = 2;
// bram[17738] = 0;
// bram[17739] = 0;
// bram[17740] = 2;
// bram[17741] = 6;
// bram[17742] = 12;
// bram[17743] = 19;
// bram[17744] = 29;
// bram[17745] = 40;
// bram[17746] = 53;
// bram[17747] = 67;
// bram[17748] = 82;
// bram[17749] = 98;
// bram[17750] = 114;
// bram[17751] = 130;
// bram[17752] = 147;
// bram[17753] = 163;
// bram[17754] = 178;
// bram[17755] = 193;
// bram[17756] = 206;
// bram[17757] = 218;
// bram[17758] = 229;
// bram[17759] = 238;
// bram[17760] = 245;
// bram[17761] = 250;
// bram[17762] = 253;
// bram[17763] = 253;
// bram[17764] = 252;
// bram[17765] = 249;
// bram[17766] = 244;
// bram[17767] = 236;
// bram[17768] = 227;
// bram[17769] = 216;
// bram[17770] = 204;
// bram[17771] = 190;
// bram[17772] = 176;
// bram[17773] = 160;
// bram[17774] = 144;
// bram[17775] = 128;
// bram[17776] = 111;
// bram[17777] = 95;
// bram[17778] = 80;
// bram[17779] = 65;
// bram[17780] = 51;
// bram[17781] = 39;
// bram[17782] = 27;
// bram[17783] = 18;
// bram[17784] = 10;
// bram[17785] = 5;
// bram[17786] = 1;
// bram[17787] = 0;
// bram[17788] = 0;
// bram[17789] = 3;
// bram[17790] = 8;
// bram[17791] = 14;
// bram[17792] = 23;
// bram[17793] = 33;
// bram[17794] = 45;
// bram[17795] = 58;
// bram[17796] = 73;
// bram[17797] = 88;
// bram[17798] = 104;
// bram[17799] = 120;
// bram[17800] = 136;
// bram[17801] = 153;
// bram[17802] = 168;
// bram[17803] = 184;
// bram[17804] = 198;
// bram[17805] = 211;
// bram[17806] = 222;
// bram[17807] = 232;
// bram[17808] = 240;
// bram[17809] = 247;
// bram[17810] = 251;
// bram[17811] = 253;
// bram[17812] = 253;
// bram[17813] = 251;
// bram[17814] = 247;
// bram[17815] = 241;
// bram[17816] = 233;
// bram[17817] = 223;
// bram[17818] = 212;
// bram[17819] = 199;
// bram[17820] = 185;
// bram[17821] = 170;
// bram[17822] = 154;
// bram[17823] = 138;
// bram[17824] = 122;
// bram[17825] = 105;
// bram[17826] = 89;
// bram[17827] = 74;
// bram[17828] = 60;
// bram[17829] = 46;
// bram[17830] = 34;
// bram[17831] = 24;
// bram[17832] = 15;
// bram[17833] = 8;
// bram[17834] = 3;
// bram[17835] = 0;
// bram[17836] = 0;
// bram[17837] = 1;
// bram[17838] = 4;
// bram[17839] = 10;
// bram[17840] = 17;
// bram[17841] = 26;
// bram[17842] = 37;
// bram[17843] = 50;
// bram[17844] = 63;
// bram[17845] = 78;
// bram[17846] = 94;
// bram[17847] = 110;
// bram[17848] = 126;
// bram[17849] = 142;
// bram[17850] = 159;
// bram[17851] = 174;
// bram[17852] = 189;
// bram[17853] = 203;
// bram[17854] = 215;
// bram[17855] = 226;
// bram[17856] = 235;
// bram[17857] = 243;
// bram[17858] = 248;
// bram[17859] = 252;
// bram[17860] = 253;
// bram[17861] = 253;
// bram[17862] = 250;
// bram[17863] = 245;
// bram[17864] = 238;
// bram[17865] = 230;
// bram[17866] = 219;
// bram[17867] = 207;
// bram[17868] = 194;
// bram[17869] = 180;
// bram[17870] = 164;
// bram[17871] = 148;
// bram[17872] = 132;
// bram[17873] = 116;
// bram[17874] = 99;
// bram[17875] = 84;
// bram[17876] = 69;
// bram[17877] = 55;
// bram[17878] = 42;
// bram[17879] = 30;
// bram[17880] = 20;
// bram[17881] = 12;
// bram[17882] = 6;
// bram[17883] = 2;
// bram[17884] = 0;
// bram[17885] = 0;
// bram[17886] = 2;
// bram[17887] = 6;
// bram[17888] = 12;
// bram[17889] = 20;
// bram[17890] = 30;
// bram[17891] = 42;
// bram[17892] = 55;
// bram[17893] = 69;
// bram[17894] = 84;
// bram[17895] = 100;
// bram[17896] = 116;
// bram[17897] = 132;
// bram[17898] = 148;
// bram[17899] = 164;
// bram[17900] = 180;
// bram[17901] = 194;
// bram[17902] = 207;
// bram[17903] = 219;
// bram[17904] = 230;
// bram[17905] = 238;
// bram[17906] = 245;
// bram[17907] = 250;
// bram[17908] = 253;
// bram[17909] = 253;
// bram[17910] = 252;
// bram[17911] = 248;
// bram[17912] = 243;
// bram[17913] = 235;
// bram[17914] = 226;
// bram[17915] = 215;
// bram[17916] = 203;
// bram[17917] = 189;
// bram[17918] = 174;
// bram[17919] = 159;
// bram[17920] = 142;
// bram[17921] = 126;
// bram[17922] = 110;
// bram[17923] = 94;
// bram[17924] = 78;
// bram[17925] = 63;
// bram[17926] = 50;
// bram[17927] = 37;
// bram[17928] = 26;
// bram[17929] = 17;
// bram[17930] = 10;
// bram[17931] = 4;
// bram[17932] = 1;
// bram[17933] = 0;
// bram[17934] = 0;
// bram[17935] = 3;
// bram[17936] = 8;
// bram[17937] = 15;
// bram[17938] = 24;
// bram[17939] = 34;
// bram[17940] = 46;
// bram[17941] = 60;
// bram[17942] = 74;
// bram[17943] = 89;
// bram[17944] = 105;
// bram[17945] = 122;
// bram[17946] = 138;
// bram[17947] = 154;
// bram[17948] = 170;
// bram[17949] = 185;
// bram[17950] = 199;
// bram[17951] = 212;
// bram[17952] = 223;
// bram[17953] = 233;
// bram[17954] = 241;
// bram[17955] = 247;
// bram[17956] = 251;
// bram[17957] = 253;
// bram[17958] = 253;
// bram[17959] = 251;
// bram[17960] = 247;
// bram[17961] = 240;
// bram[17962] = 232;
// bram[17963] = 222;
// bram[17964] = 211;
// bram[17965] = 198;
// bram[17966] = 184;
// bram[17967] = 168;
// bram[17968] = 153;
// bram[17969] = 136;
// bram[17970] = 120;
// bram[17971] = 104;
// bram[17972] = 88;
// bram[17973] = 73;
// bram[17974] = 58;
// bram[17975] = 45;
// bram[17976] = 33;
// bram[17977] = 23;
// bram[17978] = 14;
// bram[17979] = 8;
// bram[17980] = 3;
// bram[17981] = 0;
// bram[17982] = 0;
// bram[17983] = 1;
// bram[17984] = 5;
// bram[17985] = 10;
// bram[17986] = 18;
// bram[17987] = 27;
// bram[17988] = 39;
// bram[17989] = 51;
// bram[17990] = 65;
// bram[17991] = 80;
// bram[17992] = 95;
// bram[17993] = 111;
// bram[17994] = 128;
// bram[17995] = 144;
// bram[17996] = 160;
// bram[17997] = 176;
// bram[17998] = 190;
// bram[17999] = 204;
// bram[18000] = 216;
// bram[18001] = 227;
// bram[18002] = 236;
// bram[18003] = 244;
// bram[18004] = 249;
// bram[18005] = 252;
// bram[18006] = 253;
// bram[18007] = 253;
// bram[18008] = 250;
// bram[18009] = 245;
// bram[18010] = 238;
// bram[18011] = 229;
// bram[18012] = 218;
// bram[18013] = 206;
// bram[18014] = 193;
// bram[18015] = 178;
// bram[18016] = 163;
// bram[18017] = 147;
// bram[18018] = 130;
// bram[18019] = 114;
// bram[18020] = 98;
// bram[18021] = 82;
// bram[18022] = 67;
// bram[18023] = 53;
// bram[18024] = 40;
// bram[18025] = 29;
// bram[18026] = 19;
// bram[18027] = 12;
// bram[18028] = 6;
// bram[18029] = 2;
// bram[18030] = 0;
// bram[18031] = 0;
// bram[18032] = 2;
// bram[18033] = 7;
// bram[18034] = 13;
// bram[18035] = 21;
// bram[18036] = 31;
// bram[18037] = 43;
// bram[18038] = 56;
// bram[18039] = 70;
// bram[18040] = 85;
// bram[18041] = 101;
// bram[18042] = 117;
// bram[18043] = 134;
// bram[18044] = 150;
// bram[18045] = 166;
// bram[18046] = 181;
// bram[18047] = 196;
// bram[18048] = 209;
// bram[18049] = 220;
// bram[18050] = 231;
// bram[18051] = 239;
// bram[18052] = 246;
// bram[18053] = 250;
// bram[18054] = 253;
// bram[18055] = 253;
// bram[18056] = 252;
// bram[18057] = 248;
// bram[18058] = 242;
// bram[18059] = 234;
// bram[18060] = 225;
// bram[18061] = 214;
// bram[18062] = 201;
// bram[18063] = 187;
// bram[18064] = 173;
// bram[18065] = 157;
// bram[18066] = 141;
// bram[18067] = 124;
// bram[18068] = 108;
// bram[18069] = 92;
// bram[18070] = 77;
// bram[18071] = 62;
// bram[18072] = 48;
// bram[18073] = 36;
// bram[18074] = 25;
// bram[18075] = 16;
// bram[18076] = 9;
// bram[18077] = 4;
// bram[18078] = 1;
// bram[18079] = 0;
// bram[18080] = 1;
// bram[18081] = 4;
// bram[18082] = 9;
// bram[18083] = 16;
// bram[18084] = 25;
// bram[18085] = 35;
// bram[18086] = 48;
// bram[18087] = 61;
// bram[18088] = 76;
// bram[18089] = 91;
// bram[18090] = 107;
// bram[18091] = 123;
// bram[18092] = 140;
// bram[18093] = 156;
// bram[18094] = 172;
// bram[18095] = 187;
// bram[18096] = 201;
// bram[18097] = 213;
// bram[18098] = 224;
// bram[18099] = 234;
// bram[18100] = 242;
// bram[18101] = 248;
// bram[18102] = 252;
// bram[18103] = 253;
// bram[18104] = 253;
// bram[18105] = 251;
// bram[18106] = 246;
// bram[18107] = 240;
// bram[18108] = 231;
// bram[18109] = 221;
// bram[18110] = 209;
// bram[18111] = 196;
// bram[18112] = 182;
// bram[18113] = 167;
// bram[18114] = 151;
// bram[18115] = 135;
// bram[18116] = 118;
// bram[18117] = 102;
// bram[18118] = 86;
// bram[18119] = 71;
// bram[18120] = 57;
// bram[18121] = 44;
// bram[18122] = 32;
// bram[18123] = 22;
// bram[18124] = 13;
// bram[18125] = 7;
// bram[18126] = 2;
// bram[18127] = 0;
// bram[18128] = 0;
// bram[18129] = 1;
// bram[18130] = 5;
// bram[18131] = 11;
// bram[18132] = 19;
// bram[18133] = 29;
// bram[18134] = 40;
// bram[18135] = 52;
// bram[18136] = 66;
// bram[18137] = 81;
// bram[18138] = 97;
// bram[18139] = 113;
// bram[18140] = 129;
// bram[18141] = 146;
// bram[18142] = 162;
// bram[18143] = 177;
// bram[18144] = 192;
// bram[18145] = 205;
// bram[18146] = 217;
// bram[18147] = 228;
// bram[18148] = 237;
// bram[18149] = 244;
// bram[18150] = 249;
// bram[18151] = 252;
// bram[18152] = 253;
// bram[18153] = 252;
// bram[18154] = 249;
// bram[18155] = 244;
// bram[18156] = 237;
// bram[18157] = 228;
// bram[18158] = 217;
// bram[18159] = 205;
// bram[18160] = 191;
// bram[18161] = 177;
// bram[18162] = 161;
// bram[18163] = 145;
// bram[18164] = 129;
// bram[18165] = 112;
// bram[18166] = 96;
// bram[18167] = 81;
// bram[18168] = 66;
// bram[18169] = 52;
// bram[18170] = 39;
// bram[18171] = 28;
// bram[18172] = 19;
// bram[18173] = 11;
// bram[18174] = 5;
// bram[18175] = 1;
// bram[18176] = 0;
// bram[18177] = 0;
// bram[18178] = 3;
// bram[18179] = 7;
// bram[18180] = 14;
// bram[18181] = 22;
// bram[18182] = 32;
// bram[18183] = 44;
// bram[18184] = 57;
// bram[18185] = 72;
// bram[18186] = 87;
// bram[18187] = 103;
// bram[18188] = 119;
// bram[18189] = 136;
// bram[18190] = 152;
// bram[18191] = 168;
// bram[18192] = 183;
// bram[18193] = 197;
// bram[18194] = 210;
// bram[18195] = 222;
// bram[18196] = 232;
// bram[18197] = 240;
// bram[18198] = 246;
// bram[18199] = 251;
// bram[18200] = 253;
// bram[18201] = 253;
// bram[18202] = 251;
// bram[18203] = 247;
// bram[18204] = 241;
// bram[18205] = 234;
// bram[18206] = 224;
// bram[18207] = 213;
// bram[18208] = 200;
// bram[18209] = 186;
// bram[18210] = 171;
// bram[18211] = 155;
// bram[18212] = 139;
// bram[18213] = 123;
// bram[18214] = 106;
// bram[18215] = 90;
// bram[18216] = 75;
// bram[18217] = 60;
// bram[18218] = 47;
// bram[18219] = 35;
// bram[18220] = 24;
// bram[18221] = 15;
// bram[18222] = 8;
// bram[18223] = 3;
// bram[18224] = 0;
// bram[18225] = 0;
// bram[18226] = 1;
// bram[18227] = 4;
// bram[18228] = 9;
// bram[18229] = 17;
// bram[18230] = 26;
// bram[18231] = 37;
// bram[18232] = 49;
// bram[18233] = 63;
// bram[18234] = 77;
// bram[18235] = 93;
// bram[18236] = 109;
// bram[18237] = 125;
// bram[18238] = 142;
// bram[18239] = 158;
// bram[18240] = 173;
// bram[18241] = 188;
// bram[18242] = 202;
// bram[18243] = 214;
// bram[18244] = 225;
// bram[18245] = 235;
// bram[18246] = 243;
// bram[18247] = 248;
// bram[18248] = 252;
// bram[18249] = 253;
// bram[18250] = 253;
// bram[18251] = 250;
// bram[18252] = 246;
// bram[18253] = 239;
// bram[18254] = 230;
// bram[18255] = 220;
// bram[18256] = 208;
// bram[18257] = 195;
// bram[18258] = 180;
// bram[18259] = 165;
// bram[18260] = 149;
// bram[18261] = 133;
// bram[18262] = 117;
// bram[18263] = 100;
// bram[18264] = 85;
// bram[18265] = 70;
// bram[18266] = 55;
// bram[18267] = 42;
// bram[18268] = 31;
// bram[18269] = 21;
// bram[18270] = 13;
// bram[18271] = 6;
// bram[18272] = 2;
// bram[18273] = 0;
// bram[18274] = 0;
// bram[18275] = 2;
// bram[18276] = 6;
// bram[18277] = 12;
// bram[18278] = 20;
// bram[18279] = 30;
// bram[18280] = 41;
// bram[18281] = 54;
// bram[18282] = 68;
// bram[18283] = 83;
// bram[18284] = 99;
// bram[18285] = 115;
// bram[18286] = 131;
// bram[18287] = 147;
// bram[18288] = 163;
// bram[18289] = 179;
// bram[18290] = 193;
// bram[18291] = 207;
// bram[18292] = 219;
// bram[18293] = 229;
// bram[18294] = 238;
// bram[18295] = 245;
// bram[18296] = 250;
// bram[18297] = 253;
// bram[18298] = 253;
// bram[18299] = 252;
// bram[18300] = 249;
// bram[18301] = 243;
// bram[18302] = 236;
// bram[18303] = 227;
// bram[18304] = 216;
// bram[18305] = 203;
// bram[18306] = 190;
// bram[18307] = 175;
// bram[18308] = 159;
// bram[18309] = 143;
// bram[18310] = 127;
// bram[18311] = 111;
// bram[18312] = 95;
// bram[18313] = 79;
// bram[18314] = 64;
// bram[18315] = 50;
// bram[18316] = 38;
// bram[18317] = 27;
// bram[18318] = 18;
// bram[18319] = 10;
// bram[18320] = 5;
// bram[18321] = 1;
// bram[18322] = 0;
// bram[18323] = 0;
// bram[18324] = 3;
// bram[18325] = 8;
// bram[18326] = 15;
// bram[18327] = 23;
// bram[18328] = 34;
// bram[18329] = 46;
// bram[18330] = 59;
// bram[18331] = 73;
// bram[18332] = 89;
// bram[18333] = 105;
// bram[18334] = 121;
// bram[18335] = 137;
// bram[18336] = 153;
// bram[18337] = 169;
// bram[18338] = 184;
// bram[18339] = 198;
// bram[18340] = 211;
// bram[18341] = 223;
// bram[18342] = 233;
// bram[18343] = 241;
// bram[18344] = 247;
// bram[18345] = 251;
// bram[18346] = 253;
// bram[18347] = 253;
// bram[18348] = 251;
// bram[18349] = 247;
// bram[18350] = 241;
// bram[18351] = 233;
// bram[18352] = 223;
// bram[18353] = 211;
// bram[18354] = 198;
// bram[18355] = 184;
// bram[18356] = 169;
// bram[18357] = 154;
// bram[18358] = 137;
// bram[18359] = 121;
// bram[18360] = 105;
// bram[18361] = 89;
// bram[18362] = 73;
// bram[18363] = 59;
// bram[18364] = 46;
// bram[18365] = 34;
// bram[18366] = 23;
// bram[18367] = 15;
// bram[18368] = 8;
// bram[18369] = 3;
// bram[18370] = 0;
// bram[18371] = 0;
// bram[18372] = 1;
// bram[18373] = 5;
// bram[18374] = 10;
// bram[18375] = 18;
// bram[18376] = 27;
// bram[18377] = 38;
// bram[18378] = 50;
// bram[18379] = 64;
// bram[18380] = 79;
// bram[18381] = 94;
// bram[18382] = 110;
// bram[18383] = 127;
// bram[18384] = 143;
// bram[18385] = 159;
// bram[18386] = 175;
// bram[18387] = 190;
// bram[18388] = 203;
// bram[18389] = 216;
// bram[18390] = 227;
// bram[18391] = 236;
// bram[18392] = 243;
// bram[18393] = 249;
// bram[18394] = 252;
// bram[18395] = 253;
// bram[18396] = 253;
// bram[18397] = 250;
// bram[18398] = 245;
// bram[18399] = 238;
// bram[18400] = 229;
// bram[18401] = 219;
// bram[18402] = 207;
// bram[18403] = 193;
// bram[18404] = 179;
// bram[18405] = 164;
// bram[18406] = 148;
// bram[18407] = 131;
// bram[18408] = 115;
// bram[18409] = 99;
// bram[18410] = 83;
// bram[18411] = 68;
// bram[18412] = 54;
// bram[18413] = 41;
// bram[18414] = 30;
// bram[18415] = 20;
// bram[18416] = 12;
// bram[18417] = 6;
// bram[18418] = 2;
// bram[18419] = 0;
// bram[18420] = 0;
// bram[18421] = 2;
// bram[18422] = 6;
// bram[18423] = 13;
// bram[18424] = 21;
// bram[18425] = 31;
// bram[18426] = 42;
// bram[18427] = 55;
// bram[18428] = 69;
// bram[18429] = 84;
// bram[18430] = 100;
// bram[18431] = 116;
// bram[18432] = 133;
// bram[18433] = 149;
// bram[18434] = 165;
// bram[18435] = 180;
// bram[18436] = 195;
// bram[18437] = 208;
// bram[18438] = 220;
// bram[18439] = 230;
// bram[18440] = 239;
// bram[18441] = 245;
// bram[18442] = 250;
// bram[18443] = 253;
// bram[18444] = 253;
// bram[18445] = 252;
// bram[18446] = 248;
// bram[18447] = 243;
// bram[18448] = 235;
// bram[18449] = 226;
// bram[18450] = 215;
// bram[18451] = 202;
// bram[18452] = 188;
// bram[18453] = 173;
// bram[18454] = 158;
// bram[18455] = 142;
// bram[18456] = 125;
// bram[18457] = 109;
// bram[18458] = 93;
// bram[18459] = 77;
// bram[18460] = 63;
// bram[18461] = 49;
// bram[18462] = 37;
// bram[18463] = 26;
// bram[18464] = 17;
// bram[18465] = 9;
// bram[18466] = 4;
// bram[18467] = 1;
// bram[18468] = 0;
// bram[18469] = 0;
// bram[18470] = 3;
// bram[18471] = 8;
// bram[18472] = 15;
// bram[18473] = 24;
// bram[18474] = 35;
// bram[18475] = 47;
// bram[18476] = 60;
// bram[18477] = 75;
// bram[18478] = 90;
// bram[18479] = 106;
// bram[18480] = 123;
// bram[18481] = 139;
// bram[18482] = 155;
// bram[18483] = 171;
// bram[18484] = 186;
// bram[18485] = 200;
// bram[18486] = 212;
// bram[18487] = 224;
// bram[18488] = 234;
// bram[18489] = 241;
// bram[18490] = 247;
// bram[18491] = 251;
// bram[18492] = 253;
// bram[18493] = 253;
// bram[18494] = 251;
// bram[18495] = 246;
// bram[18496] = 240;
// bram[18497] = 232;
// bram[18498] = 222;
// bram[18499] = 210;
// bram[18500] = 197;
// bram[18501] = 183;
// bram[18502] = 168;
// bram[18503] = 152;
// bram[18504] = 136;
// bram[18505] = 119;
// bram[18506] = 103;
// bram[18507] = 87;
// bram[18508] = 72;
// bram[18509] = 58;
// bram[18510] = 44;
// bram[18511] = 33;
// bram[18512] = 22;
// bram[18513] = 14;
// bram[18514] = 7;
// bram[18515] = 3;
// bram[18516] = 0;
// bram[18517] = 0;
// bram[18518] = 1;
// bram[18519] = 5;
// bram[18520] = 11;
// bram[18521] = 18;
// bram[18522] = 28;
// bram[18523] = 39;
// bram[18524] = 52;
// bram[18525] = 66;
// bram[18526] = 80;
// bram[18527] = 96;
// bram[18528] = 112;
// bram[18529] = 129;
// bram[18530] = 145;
// bram[18531] = 161;
// bram[18532] = 176;
// bram[18533] = 191;
// bram[18534] = 205;
// bram[18535] = 217;
// bram[18536] = 228;
// bram[18537] = 237;
// bram[18538] = 244;
// bram[18539] = 249;
// bram[18540] = 252;
// bram[18541] = 253;
// bram[18542] = 253;
// bram[18543] = 249;
// bram[18544] = 244;
// bram[18545] = 237;
// bram[18546] = 228;
// bram[18547] = 218;
// bram[18548] = 205;
// bram[18549] = 192;
// bram[18550] = 177;
// bram[18551] = 162;
// bram[18552] = 146;
// bram[18553] = 130;
// bram[18554] = 113;
// bram[18555] = 97;
// bram[18556] = 81;
// bram[18557] = 67;
// bram[18558] = 53;
// bram[18559] = 40;
// bram[18560] = 29;
// bram[18561] = 19;
// bram[18562] = 11;
// bram[18563] = 5;
// bram[18564] = 1;
// bram[18565] = 0;
// bram[18566] = 0;
// bram[18567] = 2;
// bram[18568] = 7;
// bram[18569] = 13;
// bram[18570] = 22;
// bram[18571] = 32;
// bram[18572] = 44;
// bram[18573] = 57;
// bram[18574] = 71;
// bram[18575] = 86;
// bram[18576] = 102;
// bram[18577] = 118;
// bram[18578] = 135;
// bram[18579] = 151;
// bram[18580] = 167;
// bram[18581] = 182;
// bram[18582] = 196;
// bram[18583] = 209;
// bram[18584] = 221;
// bram[18585] = 231;
// bram[18586] = 240;
// bram[18587] = 246;
// bram[18588] = 251;
// bram[18589] = 253;
// bram[18590] = 253;
// bram[18591] = 252;
// bram[18592] = 248;
// bram[18593] = 242;
// bram[18594] = 234;
// bram[18595] = 225;
// bram[18596] = 213;
// bram[18597] = 201;
// bram[18598] = 187;
// bram[18599] = 172;
// bram[18600] = 156;
// bram[18601] = 140;
// bram[18602] = 124;
// bram[18603] = 107;
// bram[18604] = 91;
// bram[18605] = 76;
// bram[18606] = 61;
// bram[18607] = 48;
// bram[18608] = 36;
// bram[18609] = 25;
// bram[18610] = 16;
// bram[18611] = 9;
// bram[18612] = 4;
// bram[18613] = 1;
// bram[18614] = 0;
// bram[18615] = 1;
// bram[18616] = 4;
// bram[18617] = 9;
// bram[18618] = 16;
// bram[18619] = 25;
// bram[18620] = 36;
// bram[18621] = 48;
// bram[18622] = 62;
// bram[18623] = 76;
// bram[18624] = 92;
// bram[18625] = 108;
// bram[18626] = 124;
// bram[18627] = 141;
// bram[18628] = 157;
// bram[18629] = 172;
// bram[18630] = 187;
// bram[18631] = 201;
// bram[18632] = 214;
// bram[18633] = 225;
// bram[18634] = 234;
// bram[18635] = 242;
// bram[18636] = 248;
// bram[18637] = 252;
// bram[18638] = 253;
// bram[18639] = 253;
// bram[18640] = 250;
// bram[18641] = 246;
// bram[18642] = 239;
// bram[18643] = 231;
// bram[18644] = 221;
// bram[18645] = 209;
// bram[18646] = 196;
// bram[18647] = 181;
// bram[18648] = 166;
// bram[18649] = 150;
// bram[18650] = 134;
// bram[18651] = 118;
// bram[18652] = 101;
// bram[18653] = 86;
// bram[18654] = 70;
// bram[18655] = 56;
// bram[18656] = 43;
// bram[18657] = 31;
// bram[18658] = 21;
// bram[18659] = 13;
// bram[18660] = 7;
// bram[18661] = 2;
// bram[18662] = 0;
// bram[18663] = 0;
// bram[18664] = 2;
// bram[18665] = 5;
// bram[18666] = 11;
// bram[18667] = 19;
// bram[18668] = 29;
// bram[18669] = 40;
// bram[18670] = 53;
// bram[18671] = 67;
// bram[18672] = 82;
// bram[18673] = 98;
// bram[18674] = 114;
// bram[18675] = 130;
// bram[18676] = 147;
// bram[18677] = 163;
// bram[18678] = 178;
// bram[18679] = 192;
// bram[18680] = 206;
// bram[18681] = 218;
// bram[18682] = 229;
// bram[18683] = 237;
// bram[18684] = 245;
// bram[18685] = 250;
// bram[18686] = 253;
// bram[18687] = 253;
// bram[18688] = 252;
// bram[18689] = 249;
// bram[18690] = 244;
// bram[18691] = 236;
// bram[18692] = 227;
// bram[18693] = 216;
// bram[18694] = 204;
// bram[18695] = 191;
// bram[18696] = 176;
// bram[18697] = 160;
// bram[18698] = 144;
// bram[18699] = 128;
// bram[18700] = 112;
// bram[18701] = 95;
// bram[18702] = 80;
// bram[18703] = 65;
// bram[18704] = 51;
// bram[18705] = 39;
// bram[18706] = 28;
// bram[18707] = 18;
// bram[18708] = 11;
// bram[18709] = 5;
// bram[18710] = 1;
// bram[18711] = 0;
// bram[18712] = 0;
// bram[18713] = 3;
// bram[18714] = 7;
// bram[18715] = 14;
// bram[18716] = 23;
// bram[18717] = 33;
// bram[18718] = 45;
// bram[18719] = 58;
// bram[18720] = 72;
// bram[18721] = 88;
// bram[18722] = 104;
// bram[18723] = 120;
// bram[18724] = 136;
// bram[18725] = 152;
// bram[18726] = 168;
// bram[18727] = 183;
// bram[18728] = 198;
// bram[18729] = 211;
// bram[18730] = 222;
// bram[18731] = 232;
// bram[18732] = 240;
// bram[18733] = 247;
// bram[18734] = 251;
// bram[18735] = 253;
// bram[18736] = 253;
// bram[18737] = 251;
// bram[18738] = 247;
// bram[18739] = 241;
// bram[18740] = 233;
// bram[18741] = 223;
// bram[18742] = 212;
// bram[18743] = 199;
// bram[18744] = 185;
// bram[18745] = 170;
// bram[18746] = 154;
// bram[18747] = 138;
// bram[18748] = 122;
// bram[18749] = 106;
// bram[18750] = 90;
// bram[18751] = 74;
// bram[18752] = 60;
// bram[18753] = 46;
// bram[18754] = 34;
// bram[18755] = 24;
// bram[18756] = 15;
// bram[18757] = 8;
// bram[18758] = 3;
// bram[18759] = 0;
// bram[18760] = 0;
// bram[18761] = 1;
// bram[18762] = 4;
// bram[18763] = 10;
// bram[18764] = 17;
// bram[18765] = 26;
// bram[18766] = 37;
// bram[18767] = 50;
// bram[18768] = 63;
// bram[18769] = 78;
// bram[18770] = 93;
// bram[18771] = 110;
// bram[18772] = 126;
// bram[18773] = 142;
// bram[18774] = 158;
// bram[18775] = 174;
// bram[18776] = 189;
// bram[18777] = 202;
// bram[18778] = 215;
// bram[18779] = 226;
// bram[18780] = 235;
// bram[18781] = 243;
// bram[18782] = 248;
// bram[18783] = 252;
// bram[18784] = 253;
// bram[18785] = 253;
// bram[18786] = 250;
// bram[18787] = 245;
// bram[18788] = 238;
// bram[18789] = 230;
// bram[18790] = 219;
// bram[18791] = 207;
// bram[18792] = 194;
// bram[18793] = 180;
// bram[18794] = 165;
// bram[18795] = 149;
// bram[18796] = 132;
// bram[18797] = 116;
// bram[18798] = 100;
// bram[18799] = 84;
// bram[18800] = 69;
// bram[18801] = 55;
// bram[18802] = 42;
// bram[18803] = 30;
// bram[18804] = 20;
// bram[18805] = 12;
// bram[18806] = 6;
// bram[18807] = 2;
// bram[18808] = 0;
// bram[18809] = 0;
// bram[18810] = 2;
// bram[18811] = 6;
// bram[18812] = 12;
// bram[18813] = 20;
// bram[18814] = 30;
// bram[18815] = 42;
// bram[18816] = 54;
// bram[18817] = 69;
// bram[18818] = 84;
// bram[18819] = 99;
// bram[18820] = 116;
// bram[18821] = 132;
// bram[18822] = 148;
// bram[18823] = 164;
// bram[18824] = 179;
// bram[18825] = 194;
// bram[18826] = 207;
// bram[18827] = 219;
// bram[18828] = 230;
// bram[18829] = 238;
// bram[18830] = 245;
// bram[18831] = 250;
// bram[18832] = 253;
// bram[18833] = 253;
// bram[18834] = 252;
// bram[18835] = 249;
// bram[18836] = 243;
// bram[18837] = 235;
// bram[18838] = 226;
// bram[18839] = 215;
// bram[18840] = 203;
// bram[18841] = 189;
// bram[18842] = 174;
// bram[18843] = 159;
// bram[18844] = 143;
// bram[18845] = 126;
// bram[18846] = 110;
// bram[18847] = 94;
// bram[18848] = 78;
// bram[18849] = 64;
// bram[18850] = 50;
// bram[18851] = 37;
// bram[18852] = 27;
// bram[18853] = 17;
// bram[18854] = 10;
// bram[18855] = 4;
// bram[18856] = 1;
// bram[18857] = 0;
// bram[18858] = 0;
// bram[18859] = 3;
// bram[18860] = 8;
// bram[18861] = 15;
// bram[18862] = 24;
// bram[18863] = 34;
// bram[18864] = 46;
// bram[18865] = 60;
// bram[18866] = 74;
// bram[18867] = 89;
// bram[18868] = 105;
// bram[18869] = 122;
// bram[18870] = 138;
// bram[18871] = 154;
// bram[18872] = 170;
// bram[18873] = 185;
// bram[18874] = 199;
// bram[18875] = 212;
// bram[18876] = 223;
// bram[18877] = 233;
// bram[18878] = 241;
// bram[18879] = 247;
// bram[18880] = 251;
// bram[18881] = 253;
// bram[18882] = 253;
// bram[18883] = 251;
// bram[18884] = 247;
// bram[18885] = 240;
// bram[18886] = 232;
// bram[18887] = 222;
// bram[18888] = 211;
// bram[18889] = 198;
// bram[18890] = 184;
// bram[18891] = 169;
// bram[18892] = 153;
// bram[18893] = 137;
// bram[18894] = 120;
// bram[18895] = 104;
// bram[18896] = 88;
// bram[18897] = 73;
// bram[18898] = 58;
// bram[18899] = 45;
// bram[18900] = 33;
// bram[18901] = 23;
// bram[18902] = 14;
// bram[18903] = 8;
// bram[18904] = 3;
// bram[18905] = 0;
// bram[18906] = 0;
// bram[18907] = 1;
// bram[18908] = 5;
// bram[18909] = 10;
// bram[18910] = 18;
// bram[18911] = 27;
// bram[18912] = 38;
// bram[18913] = 51;
// bram[18914] = 65;
// bram[18915] = 80;
// bram[18916] = 95;
// bram[18917] = 111;
// bram[18918] = 128;
// bram[18919] = 144;
// bram[18920] = 160;
// bram[18921] = 176;
// bram[18922] = 190;
// bram[18923] = 204;
// bram[18924] = 216;
// bram[18925] = 227;
// bram[18926] = 236;
// bram[18927] = 244;
// bram[18928] = 249;
// bram[18929] = 252;
// bram[18930] = 253;
// bram[18931] = 253;
// bram[18932] = 250;
// bram[18933] = 245;
// bram[18934] = 238;
// bram[18935] = 229;
// bram[18936] = 218;
// bram[18937] = 206;
// bram[18938] = 193;
// bram[18939] = 178;
// bram[18940] = 163;
// bram[18941] = 147;
// bram[18942] = 131;
// bram[18943] = 114;
// bram[18944] = 98;
// bram[18945] = 82;
// bram[18946] = 67;
// bram[18947] = 53;
// bram[18948] = 41;
// bram[18949] = 29;
// bram[18950] = 20;
// bram[18951] = 12;
// bram[18952] = 6;
// bram[18953] = 2;
// bram[18954] = 0;
// bram[18955] = 0;
// bram[18956] = 2;
// bram[18957] = 7;
// bram[18958] = 13;
// bram[18959] = 21;
// bram[18960] = 31;
// bram[18961] = 43;
// bram[18962] = 56;
// bram[18963] = 70;
// bram[18964] = 85;
// bram[18965] = 101;
// bram[18966] = 117;
// bram[18967] = 134;
// bram[18968] = 150;
// bram[18969] = 166;
// bram[18970] = 181;
// bram[18971] = 195;
// bram[18972] = 209;
// bram[18973] = 220;
// bram[18974] = 231;
// bram[18975] = 239;
// bram[18976] = 246;
// bram[18977] = 250;
// bram[18978] = 253;
// bram[18979] = 253;
// bram[18980] = 252;
// bram[18981] = 248;
// bram[18982] = 242;
// bram[18983] = 235;
// bram[18984] = 225;
// bram[18985] = 214;
// bram[18986] = 201;
// bram[18987] = 188;
// bram[18988] = 173;
// bram[18989] = 157;
// bram[18990] = 141;
// bram[18991] = 125;
// bram[18992] = 108;
// bram[18993] = 92;
// bram[18994] = 77;
// bram[18995] = 62;
// bram[18996] = 49;
// bram[18997] = 36;
// bram[18998] = 25;
// bram[18999] = 16;
// bram[19000] = 9;
// bram[19001] = 4;
// bram[19002] = 1;
// bram[19003] = 0;
// bram[19004] = 0;
// bram[19005] = 4;
// bram[19006] = 9;
// bram[19007] = 16;
// bram[19008] = 25;
// bram[19009] = 35;
// bram[19010] = 47;
// bram[19011] = 61;
// bram[19012] = 76;
// bram[19013] = 91;
// bram[19014] = 107;
// bram[19015] = 123;
// bram[19016] = 140;
// bram[19017] = 156;
// bram[19018] = 171;
// bram[19019] = 186;
// bram[19020] = 200;
// bram[19021] = 213;
// bram[19022] = 224;
// bram[19023] = 234;
// bram[19024] = 242;
// bram[19025] = 248;
// bram[19026] = 252;
// bram[19027] = 253;
// bram[19028] = 253;
// bram[19029] = 251;
// bram[19030] = 246;
// bram[19031] = 240;
// bram[19032] = 231;
// bram[19033] = 221;
// bram[19034] = 210;
// bram[19035] = 196;
// bram[19036] = 182;
// bram[19037] = 167;
// bram[19038] = 151;
// bram[19039] = 135;
// bram[19040] = 119;
// bram[19041] = 102;
// bram[19042] = 86;
// bram[19043] = 71;
// bram[19044] = 57;
// bram[19045] = 44;
// bram[19046] = 32;
// bram[19047] = 22;
// bram[19048] = 14;
// bram[19049] = 7;
// bram[19050] = 2;
// bram[19051] = 0;
// bram[19052] = 0;
// bram[19053] = 1;
// bram[19054] = 5;
// bram[19055] = 11;
// bram[19056] = 19;
// bram[19057] = 28;
// bram[19058] = 40;
// bram[19059] = 52;
// bram[19060] = 66;
// bram[19061] = 81;
// bram[19062] = 97;
// bram[19063] = 113;
// bram[19064] = 129;
// bram[19065] = 146;
// bram[19066] = 162;
// bram[19067] = 177;
// bram[19068] = 192;
// bram[19069] = 205;
// bram[19070] = 217;
// bram[19071] = 228;
// bram[19072] = 237;
// bram[19073] = 244;
// bram[19074] = 249;
// bram[19075] = 252;
// bram[19076] = 253;
// bram[19077] = 252;
// bram[19078] = 249;
// bram[19079] = 244;
// bram[19080] = 237;
// bram[19081] = 228;
// bram[19082] = 217;
// bram[19083] = 205;
// bram[19084] = 191;
// bram[19085] = 177;
// bram[19086] = 161;
// bram[19087] = 145;
// bram[19088] = 129;
// bram[19089] = 113;
// bram[19090] = 96;
// bram[19091] = 81;
// bram[19092] = 66;
// bram[19093] = 52;
// bram[19094] = 39;
// bram[19095] = 28;
// bram[19096] = 19;
// bram[19097] = 11;
// bram[19098] = 5;
// bram[19099] = 1;
// bram[19100] = 0;
// bram[19101] = 0;
// bram[19102] = 3;
// bram[19103] = 7;
// bram[19104] = 14;
// bram[19105] = 22;
// bram[19106] = 32;
// bram[19107] = 44;
// bram[19108] = 57;
// bram[19109] = 72;
// bram[19110] = 87;
// bram[19111] = 103;
// bram[19112] = 119;
// bram[19113] = 135;
// bram[19114] = 152;
// bram[19115] = 167;
// bram[19116] = 183;
// bram[19117] = 197;
// bram[19118] = 210;
// bram[19119] = 221;
// bram[19120] = 232;
// bram[19121] = 240;
// bram[19122] = 246;
// bram[19123] = 251;
// bram[19124] = 253;
// bram[19125] = 253;
// bram[19126] = 251;
// bram[19127] = 248;
// bram[19128] = 242;
// bram[19129] = 234;
// bram[19130] = 224;
// bram[19131] = 213;
// bram[19132] = 200;
// bram[19133] = 186;
// bram[19134] = 171;
// bram[19135] = 155;
// bram[19136] = 139;
// bram[19137] = 123;
// bram[19138] = 107;
// bram[19139] = 91;
// bram[19140] = 75;
// bram[19141] = 61;
// bram[19142] = 47;
// bram[19143] = 35;
// bram[19144] = 24;
// bram[19145] = 16;
// bram[19146] = 9;
// bram[19147] = 3;
// bram[19148] = 0;
// bram[19149] = 0;
// bram[19150] = 1;
// bram[19151] = 4;
// bram[19152] = 9;
// bram[19153] = 17;
// bram[19154] = 26;
// bram[19155] = 37;
// bram[19156] = 49;
// bram[19157] = 62;
// bram[19158] = 77;
// bram[19159] = 93;
// bram[19160] = 109;
// bram[19161] = 125;
// bram[19162] = 141;
// bram[19163] = 157;
// bram[19164] = 173;
// bram[19165] = 188;
// bram[19166] = 202;
// bram[19167] = 214;
// bram[19168] = 225;
// bram[19169] = 235;
// bram[19170] = 242;
// bram[19171] = 248;
// bram[19172] = 252;
// bram[19173] = 253;
// bram[19174] = 253;
// bram[19175] = 250;
// bram[19176] = 246;
// bram[19177] = 239;
// bram[19178] = 230;
// bram[19179] = 220;
// bram[19180] = 208;
// bram[19181] = 195;
// bram[19182] = 181;
// bram[19183] = 165;
// bram[19184] = 150;
// bram[19185] = 133;
// bram[19186] = 117;
// bram[19187] = 101;
// bram[19188] = 85;
// bram[19189] = 70;
// bram[19190] = 56;
// bram[19191] = 43;
// bram[19192] = 31;
// bram[19193] = 21;
// bram[19194] = 13;
// bram[19195] = 6;
// bram[19196] = 2;
// bram[19197] = 0;
// bram[19198] = 0;
// bram[19199] = 2;
// bram[19200] = 6;
// bram[19201] = 12;
// bram[19202] = 20;
// bram[19203] = 30;
// bram[19204] = 41;
// bram[19205] = 54;
// bram[19206] = 68;
// bram[19207] = 83;
// bram[19208] = 98;
// bram[19209] = 115;
// bram[19210] = 131;
// bram[19211] = 147;
// bram[19212] = 163;
// bram[19213] = 179;
// bram[19214] = 193;
// bram[19215] = 206;
// bram[19216] = 219;
// bram[19217] = 229;
// bram[19218] = 238;
// bram[19219] = 245;
// bram[19220] = 250;
// bram[19221] = 253;
// bram[19222] = 253;
// bram[19223] = 252;
// bram[19224] = 249;
// bram[19225] = 243;
// bram[19226] = 236;
// bram[19227] = 227;
// bram[19228] = 216;
// bram[19229] = 204;
// bram[19230] = 190;
// bram[19231] = 175;
// bram[19232] = 160;
// bram[19233] = 144;
// bram[19234] = 127;
// bram[19235] = 111;
// bram[19236] = 95;
// bram[19237] = 79;
// bram[19238] = 64;
// bram[19239] = 51;
// bram[19240] = 38;
// bram[19241] = 27;
// bram[19242] = 18;
// bram[19243] = 10;
// bram[19244] = 5;
// bram[19245] = 1;
// bram[19246] = 0;
// bram[19247] = 0;
// bram[19248] = 3;
// bram[19249] = 8;
// bram[19250] = 14;
// bram[19251] = 23;
// bram[19252] = 34;
// bram[19253] = 45;
// bram[19254] = 59;
// bram[19255] = 73;
// bram[19256] = 88;
// bram[19257] = 104;
// bram[19258] = 121;
// bram[19259] = 137;
// bram[19260] = 153;
// bram[19261] = 169;
// bram[19262] = 184;
// bram[19263] = 198;
// bram[19264] = 211;
// bram[19265] = 223;
// bram[19266] = 232;
// bram[19267] = 241;
// bram[19268] = 247;
// bram[19269] = 251;
// bram[19270] = 253;
// bram[19271] = 253;
// bram[19272] = 251;
// bram[19273] = 247;
// bram[19274] = 241;
// bram[19275] = 233;
// bram[19276] = 223;
// bram[19277] = 211;
// bram[19278] = 199;
// bram[19279] = 185;
// bram[19280] = 170;
// bram[19281] = 154;
// bram[19282] = 138;
// bram[19283] = 121;
// bram[19284] = 105;
// bram[19285] = 89;
// bram[19286] = 74;
// bram[19287] = 59;
// bram[19288] = 46;
// bram[19289] = 34;
// bram[19290] = 23;
// bram[19291] = 15;
// bram[19292] = 8;
// bram[19293] = 3;
// bram[19294] = 0;
// bram[19295] = 0;
// bram[19296] = 1;
// bram[19297] = 4;
// bram[19298] = 10;
// bram[19299] = 17;
// bram[19300] = 27;
// bram[19301] = 38;
// bram[19302] = 50;
// bram[19303] = 64;
// bram[19304] = 79;
// bram[19305] = 94;
// bram[19306] = 110;
// bram[19307] = 127;
// bram[19308] = 143;
// bram[19309] = 159;
// bram[19310] = 175;
// bram[19311] = 189;
// bram[19312] = 203;
// bram[19313] = 215;
// bram[19314] = 226;
// bram[19315] = 236;
// bram[19316] = 243;
// bram[19317] = 249;
// bram[19318] = 252;
// bram[19319] = 253;
// bram[19320] = 253;
// bram[19321] = 250;
// bram[19322] = 245;
// bram[19323] = 238;
// bram[19324] = 229;
// bram[19325] = 219;
// bram[19326] = 207;
// bram[19327] = 194;
// bram[19328] = 179;
// bram[19329] = 164;
// bram[19330] = 148;
// bram[19331] = 132;
// bram[19332] = 115;
// bram[19333] = 99;
// bram[19334] = 83;
// bram[19335] = 68;
// bram[19336] = 54;
// bram[19337] = 41;
// bram[19338] = 30;
// bram[19339] = 20;
// bram[19340] = 12;
// bram[19341] = 6;
// bram[19342] = 2;
// bram[19343] = 0;
// bram[19344] = 0;
// bram[19345] = 2;
// bram[19346] = 6;
// bram[19347] = 13;
// bram[19348] = 21;
// bram[19349] = 31;
// bram[19350] = 42;
// bram[19351] = 55;
// bram[19352] = 69;
// bram[19353] = 84;
// bram[19354] = 100;
// bram[19355] = 116;
// bram[19356] = 133;
// bram[19357] = 149;
// bram[19358] = 165;
// bram[19359] = 180;
// bram[19360] = 195;
// bram[19361] = 208;
// bram[19362] = 220;
// bram[19363] = 230;
// bram[19364] = 239;
// bram[19365] = 245;
// bram[19366] = 250;
// bram[19367] = 253;
// bram[19368] = 253;
// bram[19369] = 252;
// bram[19370] = 248;
// bram[19371] = 243;
// bram[19372] = 235;
// bram[19373] = 226;
// bram[19374] = 215;
// bram[19375] = 202;
// bram[19376] = 188;
// bram[19377] = 174;
// bram[19378] = 158;
// bram[19379] = 142;
// bram[19380] = 126;
// bram[19381] = 109;
// bram[19382] = 93;
// bram[19383] = 78;
// bram[19384] = 63;
// bram[19385] = 49;
// bram[19386] = 37;
// bram[19387] = 26;
// bram[19388] = 17;
// bram[19389] = 10;
// bram[19390] = 4;
// bram[19391] = 1;
// bram[19392] = 0;
// bram[19393] = 0;
// bram[19394] = 3;
// bram[19395] = 8;
// bram[19396] = 15;
// bram[19397] = 24;
// bram[19398] = 35;
// bram[19399] = 47;
// bram[19400] = 60;
// bram[19401] = 75;
// bram[19402] = 90;
// bram[19403] = 106;
// bram[19404] = 122;
// bram[19405] = 139;
// bram[19406] = 155;
// bram[19407] = 171;
// bram[19408] = 186;
// bram[19409] = 200;
// bram[19410] = 212;
// bram[19411] = 224;
// bram[19412] = 233;
// bram[19413] = 241;
// bram[19414] = 247;
// bram[19415] = 251;
// bram[19416] = 253;
// bram[19417] = 253;
// bram[19418] = 251;
// bram[19419] = 246;
// bram[19420] = 240;
// bram[19421] = 232;
// bram[19422] = 222;
// bram[19423] = 210;
// bram[19424] = 197;
// bram[19425] = 183;
// bram[19426] = 168;
// bram[19427] = 152;
// bram[19428] = 136;
// bram[19429] = 119;
// bram[19430] = 103;
// bram[19431] = 87;
// bram[19432] = 72;
// bram[19433] = 58;
// bram[19434] = 45;
// bram[19435] = 33;
// bram[19436] = 22;
// bram[19437] = 14;
// bram[19438] = 7;
// bram[19439] = 3;
// bram[19440] = 0;
// bram[19441] = 0;
// bram[19442] = 1;
// bram[19443] = 5;
// bram[19444] = 11;
// bram[19445] = 18;
// bram[19446] = 28;
// bram[19447] = 39;
// bram[19448] = 52;
// bram[19449] = 65;
// bram[19450] = 80;
// bram[19451] = 96;
// bram[19452] = 112;
// bram[19453] = 128;
// bram[19454] = 145;
// bram[19455] = 161;
// bram[19456] = 176;
// bram[19457] = 191;
// bram[19458] = 204;
// bram[19459] = 217;
// bram[19460] = 227;
// bram[19461] = 237;
// bram[19462] = 244;
// bram[19463] = 249;
// bram[19464] = 252;
// bram[19465] = 253;
// bram[19466] = 253;
// bram[19467] = 249;
// bram[19468] = 244;
// bram[19469] = 237;
// bram[19470] = 228;
// bram[19471] = 218;
// bram[19472] = 206;
// bram[19473] = 192;
// bram[19474] = 178;
// bram[19475] = 162;
// bram[19476] = 146;
// bram[19477] = 130;
// bram[19478] = 113;
// bram[19479] = 97;
// bram[19480] = 82;
// bram[19481] = 67;
// bram[19482] = 53;
// bram[19483] = 40;
// bram[19484] = 29;
// bram[19485] = 19;
// bram[19486] = 11;
// bram[19487] = 5;
// bram[19488] = 1;
// bram[19489] = 0;
// bram[19490] = 0;
// bram[19491] = 2;
// bram[19492] = 7;
// bram[19493] = 13;
// bram[19494] = 22;
// bram[19495] = 32;
// bram[19496] = 43;
// bram[19497] = 56;
// bram[19498] = 71;
// bram[19499] = 86;
// bram[19500] = 102;
// bram[19501] = 118;
// bram[19502] = 134;
// bram[19503] = 151;
// bram[19504] = 167;
// bram[19505] = 182;
// bram[19506] = 196;
// bram[19507] = 209;
// bram[19508] = 221;
// bram[19509] = 231;
// bram[19510] = 239;
// bram[19511] = 246;
// bram[19512] = 251;
// bram[19513] = 253;
// bram[19514] = 253;
// bram[19515] = 252;
// bram[19516] = 248;
// bram[19517] = 242;
// bram[19518] = 234;
// bram[19519] = 225;
// bram[19520] = 213;
// bram[19521] = 201;
// bram[19522] = 187;
// bram[19523] = 172;
// bram[19524] = 156;
// bram[19525] = 140;
// bram[19526] = 124;
// bram[19527] = 107;
// bram[19528] = 91;
// bram[19529] = 76;
// bram[19530] = 61;
// bram[19531] = 48;
// bram[19532] = 36;
// bram[19533] = 25;
// bram[19534] = 16;
// bram[19535] = 9;
// bram[19536] = 4;
// bram[19537] = 1;
// bram[19538] = 0;
// bram[19539] = 1;
// bram[19540] = 4;
// bram[19541] = 9;
// bram[19542] = 16;
// bram[19543] = 25;
// bram[19544] = 36;
// bram[19545] = 48;
// bram[19546] = 62;
// bram[19547] = 76;
// bram[19548] = 92;
// bram[19549] = 108;
// bram[19550] = 124;
// bram[19551] = 140;
// bram[19552] = 157;
// bram[19553] = 172;
// bram[19554] = 187;
// bram[19555] = 201;
// bram[19556] = 214;
// bram[19557] = 225;
// bram[19558] = 234;
// bram[19559] = 242;
// bram[19560] = 248;
// bram[19561] = 252;
// bram[19562] = 253;
// bram[19563] = 253;
// bram[19564] = 250;
// bram[19565] = 246;
// bram[19566] = 239;
// bram[19567] = 231;
// bram[19568] = 221;
// bram[19569] = 209;
// bram[19570] = 196;
// bram[19571] = 182;
// bram[19572] = 166;
// bram[19573] = 150;
// bram[19574] = 134;
// bram[19575] = 118;
// bram[19576] = 102;
// bram[19577] = 86;
// bram[19578] = 71;
// bram[19579] = 56;
// bram[19580] = 43;
// bram[19581] = 32;
// bram[19582] = 22;
// bram[19583] = 13;
// bram[19584] = 7;
// bram[19585] = 2;
// bram[19586] = 0;
// bram[19587] = 0;
// bram[19588] = 1;
// bram[19589] = 5;
// bram[19590] = 11;
// bram[19591] = 19;
// bram[19592] = 29;
// bram[19593] = 40;
// bram[19594] = 53;
// bram[19595] = 67;
// bram[19596] = 82;
// bram[19597] = 97;
// bram[19598] = 114;
// bram[19599] = 130;
// bram[19600] = 146;
// bram[19601] = 162;
// bram[19602] = 178;
// bram[19603] = 192;
// bram[19604] = 206;
// bram[19605] = 218;
// bram[19606] = 228;
// bram[19607] = 237;
// bram[19608] = 244;
// bram[19609] = 250;
// bram[19610] = 253;
// bram[19611] = 253;
// bram[19612] = 252;
// bram[19613] = 249;
// bram[19614] = 244;
// bram[19615] = 236;
// bram[19616] = 227;
// bram[19617] = 217;
// bram[19618] = 204;
// bram[19619] = 191;
// bram[19620] = 176;
// bram[19621] = 161;
// bram[19622] = 144;
// bram[19623] = 128;
// bram[19624] = 112;
// bram[19625] = 96;
// bram[19626] = 80;
// bram[19627] = 65;
// bram[19628] = 51;
// bram[19629] = 39;
// bram[19630] = 28;
// bram[19631] = 18;
// bram[19632] = 11;
// bram[19633] = 5;
// bram[19634] = 1;
// bram[19635] = 0;
// bram[19636] = 0;
// bram[19637] = 3;
// bram[19638] = 7;
// bram[19639] = 14;
// bram[19640] = 23;
// bram[19641] = 33;
// bram[19642] = 45;
// bram[19643] = 58;
// bram[19644] = 72;
// bram[19645] = 87;
// bram[19646] = 103;
// bram[19647] = 120;
// bram[19648] = 136;
// bram[19649] = 152;
// bram[19650] = 168;
// bram[19651] = 183;
// bram[19652] = 197;
// bram[19653] = 210;
// bram[19654] = 222;
// bram[19655] = 232;
// bram[19656] = 240;
// bram[19657] = 247;
// bram[19658] = 251;
// bram[19659] = 253;
// bram[19660] = 253;
// bram[19661] = 251;
// bram[19662] = 247;
// bram[19663] = 241;
// bram[19664] = 233;
// bram[19665] = 224;
// bram[19666] = 212;
// bram[19667] = 199;
// bram[19668] = 185;
// bram[19669] = 170;
// bram[19670] = 155;
// bram[19671] = 139;
// bram[19672] = 122;
// bram[19673] = 106;
// bram[19674] = 90;
// bram[19675] = 74;
// bram[19676] = 60;
// bram[19677] = 47;
// bram[19678] = 35;
// bram[19679] = 24;
// bram[19680] = 15;
// bram[19681] = 8;
// bram[19682] = 3;
// bram[19683] = 0;
// bram[19684] = 0;
// bram[19685] = 1;
// bram[19686] = 4;
// bram[19687] = 10;
// bram[19688] = 17;
// bram[19689] = 26;
// bram[19690] = 37;
// bram[19691] = 49;
// bram[19692] = 63;
// bram[19693] = 78;
// bram[19694] = 93;
// bram[19695] = 109;
// bram[19696] = 126;
// bram[19697] = 142;
// bram[19698] = 158;
// bram[19699] = 174;
// bram[19700] = 189;
// bram[19701] = 202;
// bram[19702] = 215;
// bram[19703] = 226;
// bram[19704] = 235;
// bram[19705] = 243;
// bram[19706] = 248;
// bram[19707] = 252;
// bram[19708] = 253;
// bram[19709] = 253;
// bram[19710] = 250;
// bram[19711] = 245;
// bram[19712] = 239;
// bram[19713] = 230;
// bram[19714] = 220;
// bram[19715] = 208;
// bram[19716] = 194;
// bram[19717] = 180;
// bram[19718] = 165;
// bram[19719] = 149;
// bram[19720] = 132;
// bram[19721] = 116;
// bram[19722] = 100;
// bram[19723] = 84;
// bram[19724] = 69;
// bram[19725] = 55;
// bram[19726] = 42;
// bram[19727] = 30;
// bram[19728] = 21;
// bram[19729] = 12;
// bram[19730] = 6;
// bram[19731] = 2;
// bram[19732] = 0;
// bram[19733] = 0;
// bram[19734] = 2;
// bram[19735] = 6;
// bram[19736] = 12;
// bram[19737] = 20;
// bram[19738] = 30;
// bram[19739] = 41;
// bram[19740] = 54;
// bram[19741] = 68;
// bram[19742] = 83;
// bram[19743] = 99;
// bram[19744] = 115;
// bram[19745] = 132;
// bram[19746] = 148;
// bram[19747] = 164;
// bram[19748] = 179;
// bram[19749] = 194;
// bram[19750] = 207;
// bram[19751] = 219;
// bram[19752] = 229;
// bram[19753] = 238;
// bram[19754] = 245;
// bram[19755] = 250;
// bram[19756] = 253;
// bram[19757] = 253;
// bram[19758] = 252;
// bram[19759] = 249;
// bram[19760] = 243;
// bram[19761] = 236;
// bram[19762] = 226;
// bram[19763] = 215;
// bram[19764] = 203;
// bram[19765] = 189;
// bram[19766] = 174;
// bram[19767] = 159;
// bram[19768] = 143;
// bram[19769] = 126;
// bram[19770] = 110;
// bram[19771] = 94;
// bram[19772] = 78;
// bram[19773] = 64;
// bram[19774] = 50;
// bram[19775] = 38;
// bram[19776] = 27;
// bram[19777] = 17;
// bram[19778] = 10;
// bram[19779] = 4;
// bram[19780] = 1;
// bram[19781] = 0;
// bram[19782] = 0;
// bram[19783] = 3;
// bram[19784] = 8;
// bram[19785] = 15;
// bram[19786] = 24;
// bram[19787] = 34;
// bram[19788] = 46;
// bram[19789] = 59;
// bram[19790] = 74;
// bram[19791] = 89;
// bram[19792] = 105;
// bram[19793] = 121;
// bram[19794] = 138;
// bram[19795] = 154;
// bram[19796] = 170;
// bram[19797] = 185;
// bram[19798] = 199;
// bram[19799] = 212;
// bram[19800] = 223;
// bram[19801] = 233;
// bram[19802] = 241;
// bram[19803] = 247;
// bram[19804] = 251;
// bram[19805] = 253;
// bram[19806] = 253;
// bram[19807] = 251;
// bram[19808] = 247;
// bram[19809] = 241;
// bram[19810] = 232;
// bram[19811] = 222;
// bram[19812] = 211;
// bram[19813] = 198;
// bram[19814] = 184;
// bram[19815] = 169;
// bram[19816] = 153;
// bram[19817] = 137;
// bram[19818] = 120;
// bram[19819] = 104;
// bram[19820] = 88;
// bram[19821] = 73;
// bram[19822] = 59;
// bram[19823] = 45;
// bram[19824] = 33;
// bram[19825] = 23;
// bram[19826] = 14;
// bram[19827] = 8;
// bram[19828] = 3;
// bram[19829] = 0;
// bram[19830] = 0;
// bram[19831] = 1;
// bram[19832] = 5;
// bram[19833] = 10;
// bram[19834] = 18;
// bram[19835] = 27;
// bram[19836] = 38;
// bram[19837] = 51;
// bram[19838] = 65;
// bram[19839] = 79;
// bram[19840] = 95;
// bram[19841] = 111;
// bram[19842] = 127;
// bram[19843] = 144;
// bram[19844] = 160;
// bram[19845] = 175;
// bram[19846] = 190;
// bram[19847] = 204;
// bram[19848] = 216;
// bram[19849] = 227;
// bram[19850] = 236;
// bram[19851] = 243;
// bram[19852] = 249;
// bram[19853] = 252;
// bram[19854] = 253;
// bram[19855] = 253;
// bram[19856] = 250;
// bram[19857] = 245;
// bram[19858] = 238;
// bram[19859] = 229;
// bram[19860] = 218;
// bram[19861] = 206;
// bram[19862] = 193;
// bram[19863] = 178;
// bram[19864] = 163;
// bram[19865] = 147;
// bram[19866] = 131;
// bram[19867] = 114;
// bram[19868] = 98;
// bram[19869] = 82;
// bram[19870] = 68;
// bram[19871] = 54;
// bram[19872] = 41;
// bram[19873] = 29;
// bram[19874] = 20;
// bram[19875] = 12;
// bram[19876] = 6;
// bram[19877] = 2;
// bram[19878] = 0;
// bram[19879] = 0;
// bram[19880] = 2;
// bram[19881] = 6;
// bram[19882] = 13;
// bram[19883] = 21;
// bram[19884] = 31;
// bram[19885] = 43;
// bram[19886] = 56;
// bram[19887] = 70;
// bram[19888] = 85;
// bram[19889] = 101;
// bram[19890] = 117;
// bram[19891] = 133;
// bram[19892] = 150;
// bram[19893] = 166;
// bram[19894] = 181;
// bram[19895] = 195;
// bram[19896] = 208;
// bram[19897] = 220;
// bram[19898] = 230;
// bram[19899] = 239;
// bram[19900] = 246;
// bram[19901] = 250;
// bram[19902] = 253;
// bram[19903] = 253;
// bram[19904] = 252;
// bram[19905] = 248;
// bram[19906] = 242;
// bram[19907] = 235;
// bram[19908] = 225;
// bram[19909] = 214;
// bram[19910] = 202;
// bram[19911] = 188;
// bram[19912] = 173;
// bram[19913] = 157;
// bram[19914] = 141;
// bram[19915] = 125;
// bram[19916] = 108;
// bram[19917] = 92;
// bram[19918] = 77;
// bram[19919] = 62;
// bram[19920] = 49;
// bram[19921] = 36;
// bram[19922] = 26;
// bram[19923] = 17;
// bram[19924] = 9;
// bram[19925] = 4;
// bram[19926] = 1;
// bram[19927] = 0;
// bram[19928] = 0;
// bram[19929] = 4;
// bram[19930] = 9;
// bram[19931] = 16;
// bram[19932] = 25;
// bram[19933] = 35;
// bram[19934] = 47;
// bram[19935] = 61;
// bram[19936] = 75;
// bram[19937] = 91;
// bram[19938] = 107;
// bram[19939] = 123;
// bram[19940] = 139;
// bram[19941] = 156;
// bram[19942] = 171;
// bram[19943] = 186;
// bram[19944] = 200;
// bram[19945] = 213;
// bram[19946] = 224;
// bram[19947] = 234;
// bram[19948] = 242;
// bram[19949] = 248;
// bram[19950] = 252;
// bram[19951] = 253;
// bram[19952] = 253;
// bram[19953] = 251;
// bram[19954] = 246;
// bram[19955] = 240;
// bram[19956] = 231;
// bram[19957] = 221;
// bram[19958] = 210;
// bram[19959] = 197;
// bram[19960] = 182;
// bram[19961] = 167;
// bram[19962] = 151;
// bram[19963] = 135;
// bram[19964] = 119;
// bram[19965] = 102;
// bram[19966] = 87;
// bram[19967] = 71;
// bram[19968] = 57;
// bram[19969] = 44;
// bram[19970] = 32;
// bram[19971] = 22;
// bram[19972] = 14;
// bram[19973] = 7;
// bram[19974] = 2;
// bram[19975] = 0;
// bram[19976] = 0;
// bram[19977] = 1;
// bram[19978] = 5;
// bram[19979] = 11;
// bram[19980] = 19;
// bram[19981] = 28;
// bram[19982] = 39;
// bram[19983] = 52;
// bram[19984] = 66;
// bram[19985] = 81;
// bram[19986] = 97;
// bram[19987] = 113;
// bram[19988] = 129;
// bram[19989] = 145;
// bram[19990] = 161;
// bram[19991] = 177;
// bram[19992] = 191;
// bram[19993] = 205;
// bram[19994] = 217;
// bram[19995] = 228;
// bram[19996] = 237;
// bram[19997] = 244;
// bram[19998] = 249;
// bram[19999] = 252;
// bram[20000] = 254;
// bram[20001] = 252;
// bram[20002] = 249;
// bram[20003] = 244;
// bram[20004] = 237;
// bram[20005] = 228;
// bram[20006] = 217;
// bram[20007] = 205;
// bram[20008] = 191;
// bram[20009] = 177;
// bram[20010] = 161;
// bram[20011] = 145;
// bram[20012] = 129;
// bram[20013] = 113;
// bram[20014] = 97;
// bram[20015] = 81;
// bram[20016] = 66;
// bram[20017] = 52;
// bram[20018] = 39;
// bram[20019] = 28;
// bram[20020] = 19;
// bram[20021] = 11;
// bram[20022] = 5;
// bram[20023] = 1;
// bram[20024] = 0;
// bram[20025] = 0;
// bram[20026] = 2;
// bram[20027] = 7;
// bram[20028] = 14;
// bram[20029] = 22;
// bram[20030] = 32;
// bram[20031] = 44;
// bram[20032] = 57;
// bram[20033] = 71;
// bram[20034] = 87;
// bram[20035] = 102;
// bram[20036] = 119;
// bram[20037] = 135;
// bram[20038] = 151;
// bram[20039] = 167;
// bram[20040] = 182;
// bram[20041] = 197;
// bram[20042] = 210;
// bram[20043] = 221;
// bram[20044] = 231;
// bram[20045] = 240;
// bram[20046] = 246;
// bram[20047] = 251;
// bram[20048] = 253;
// bram[20049] = 253;
// bram[20050] = 252;
// bram[20051] = 248;
// bram[20052] = 242;
// bram[20053] = 234;
// bram[20054] = 224;
// bram[20055] = 213;
// bram[20056] = 200;
// bram[20057] = 186;
// bram[20058] = 171;
// bram[20059] = 156;
// bram[20060] = 139;
// bram[20061] = 123;
// bram[20062] = 107;
// bram[20063] = 91;
// bram[20064] = 75;
// bram[20065] = 61;
// bram[20066] = 47;
// bram[20067] = 35;
// bram[20068] = 25;
// bram[20069] = 16;
// bram[20070] = 9;
// bram[20071] = 4;
// bram[20072] = 0;
// bram[20073] = 0;
// bram[20074] = 1;
// bram[20075] = 4;
// bram[20076] = 9;
// bram[20077] = 17;
// bram[20078] = 26;
// bram[20079] = 36;
// bram[20080] = 49;
// bram[20081] = 62;
// bram[20082] = 77;
// bram[20083] = 92;
// bram[20084] = 108;
// bram[20085] = 125;
// bram[20086] = 141;
// bram[20087] = 157;
// bram[20088] = 173;
// bram[20089] = 188;
// bram[20090] = 202;
// bram[20091] = 214;
// bram[20092] = 225;
// bram[20093] = 235;
// bram[20094] = 242;
// bram[20095] = 248;
// bram[20096] = 252;
// bram[20097] = 253;
// bram[20098] = 253;
// bram[20099] = 250;
// bram[20100] = 246;
// bram[20101] = 239;
// bram[20102] = 230;
// bram[20103] = 220;
// bram[20104] = 208;
// bram[20105] = 195;
// bram[20106] = 181;
// bram[20107] = 166;
// bram[20108] = 150;
// bram[20109] = 133;
// bram[20110] = 117;
// bram[20111] = 101;
// bram[20112] = 85;
// bram[20113] = 70;
// bram[20114] = 56;
// bram[20115] = 43;
// bram[20116] = 31;
// bram[20117] = 21;
// bram[20118] = 13;
// bram[20119] = 6;
// bram[20120] = 2;
// bram[20121] = 0;
// bram[20122] = 0;
// bram[20123] = 2;
// bram[20124] = 6;
// bram[20125] = 12;
// bram[20126] = 20;
// bram[20127] = 29;
// bram[20128] = 41;
// bram[20129] = 54;
// bram[20130] = 68;
// bram[20131] = 82;
// bram[20132] = 98;
// bram[20133] = 114;
// bram[20134] = 131;
// bram[20135] = 147;
// bram[20136] = 163;
// bram[20137] = 178;
// bram[20138] = 193;
// bram[20139] = 206;
// bram[20140] = 218;
// bram[20141] = 229;
// bram[20142] = 238;
// bram[20143] = 245;
// bram[20144] = 250;
// bram[20145] = 253;
// bram[20146] = 253;
// bram[20147] = 252;
// bram[20148] = 249;
// bram[20149] = 243;
// bram[20150] = 236;
// bram[20151] = 227;
// bram[20152] = 216;
// bram[20153] = 204;
// bram[20154] = 190;
// bram[20155] = 175;
// bram[20156] = 160;
// bram[20157] = 144;
// bram[20158] = 127;
// bram[20159] = 111;
// bram[20160] = 95;
// bram[20161] = 79;
// bram[20162] = 65;
// bram[20163] = 51;
// bram[20164] = 38;
// bram[20165] = 27;
// bram[20166] = 18;
// bram[20167] = 10;
// bram[20168] = 5;
// bram[20169] = 1;
// bram[20170] = 0;
// bram[20171] = 0;
// bram[20172] = 3;
// bram[20173] = 8;
// bram[20174] = 14;
// bram[20175] = 23;
// bram[20176] = 33;
// bram[20177] = 45;
// bram[20178] = 59;
// bram[20179] = 73;
// bram[20180] = 88;
// bram[20181] = 104;
// bram[20182] = 120;
// bram[20183] = 137;
// bram[20184] = 153;
// bram[20185] = 169;
// bram[20186] = 184;
// bram[20187] = 198;
// bram[20188] = 211;
// bram[20189] = 222;
// bram[20190] = 232;
// bram[20191] = 241;
// bram[20192] = 247;
// bram[20193] = 251;
// bram[20194] = 253;
// bram[20195] = 253;
// bram[20196] = 251;
// bram[20197] = 247;
// bram[20198] = 241;
// bram[20199] = 233;
// bram[20200] = 223;
// bram[20201] = 212;
// bram[20202] = 199;
// bram[20203] = 185;
// bram[20204] = 170;
// bram[20205] = 154;
// bram[20206] = 138;
// bram[20207] = 121;
// bram[20208] = 105;
// bram[20209] = 89;
// bram[20210] = 74;
// bram[20211] = 59;
// bram[20212] = 46;
// bram[20213] = 34;
// bram[20214] = 24;
// bram[20215] = 15;
// bram[20216] = 8;
// bram[20217] = 3;
// bram[20218] = 0;
// bram[20219] = 0;
// bram[20220] = 1;
// bram[20221] = 4;
// bram[20222] = 10;
// bram[20223] = 17;
// bram[20224] = 27;
// bram[20225] = 38;
// bram[20226] = 50;
// bram[20227] = 64;
// bram[20228] = 78;
// bram[20229] = 94;
// bram[20230] = 110;
// bram[20231] = 126;
// bram[20232] = 143;
// bram[20233] = 159;
// bram[20234] = 174;
// bram[20235] = 189;
// bram[20236] = 203;
// bram[20237] = 215;
// bram[20238] = 226;
// bram[20239] = 236;
// bram[20240] = 243;
// bram[20241] = 249;
// bram[20242] = 252;
// bram[20243] = 253;
// bram[20244] = 253;
// bram[20245] = 250;
// bram[20246] = 245;
// bram[20247] = 238;
// bram[20248] = 229;
// bram[20249] = 219;
// bram[20250] = 207;
// bram[20251] = 194;
// bram[20252] = 179;
// bram[20253] = 164;
// bram[20254] = 148;
// bram[20255] = 132;
// bram[20256] = 115;
// bram[20257] = 99;
// bram[20258] = 83;
// bram[20259] = 68;
// bram[20260] = 54;
// bram[20261] = 41;
// bram[20262] = 30;
// bram[20263] = 20;
// bram[20264] = 12;
// bram[20265] = 6;
// bram[20266] = 2;
// bram[20267] = 0;
// bram[20268] = 0;
// bram[20269] = 2;
// bram[20270] = 6;
// bram[20271] = 12;
// bram[20272] = 21;
// bram[20273] = 30;
// bram[20274] = 42;
// bram[20275] = 55;
// bram[20276] = 69;
// bram[20277] = 84;
// bram[20278] = 100;
// bram[20279] = 116;
// bram[20280] = 132;
// bram[20281] = 149;
// bram[20282] = 165;
// bram[20283] = 180;
// bram[20284] = 194;
// bram[20285] = 208;
// bram[20286] = 220;
// bram[20287] = 230;
// bram[20288] = 239;
// bram[20289] = 245;
// bram[20290] = 250;
// bram[20291] = 253;
// bram[20292] = 253;
// bram[20293] = 252;
// bram[20294] = 248;
// bram[20295] = 243;
// bram[20296] = 235;
// bram[20297] = 226;
// bram[20298] = 215;
// bram[20299] = 202;
// bram[20300] = 189;
// bram[20301] = 174;
// bram[20302] = 158;
// bram[20303] = 142;
// bram[20304] = 126;
// bram[20305] = 109;
// bram[20306] = 93;
// bram[20307] = 78;
// bram[20308] = 63;
// bram[20309] = 49;
// bram[20310] = 37;
// bram[20311] = 26;
// bram[20312] = 17;
// bram[20313] = 10;
// bram[20314] = 4;
// bram[20315] = 1;
// bram[20316] = 0;
// bram[20317] = 0;
// bram[20318] = 3;
// bram[20319] = 8;
// bram[20320] = 15;
// bram[20321] = 24;
// bram[20322] = 35;
// bram[20323] = 47;
// bram[20324] = 60;
// bram[20325] = 74;
// bram[20326] = 90;
// bram[20327] = 106;
// bram[20328] = 122;
// bram[20329] = 139;
// bram[20330] = 155;
// bram[20331] = 170;
// bram[20332] = 185;
// bram[20333] = 199;
// bram[20334] = 212;
// bram[20335] = 224;
// bram[20336] = 233;
// bram[20337] = 241;
// bram[20338] = 247;
// bram[20339] = 251;
// bram[20340] = 253;
// bram[20341] = 253;
// bram[20342] = 251;
// bram[20343] = 247;
// bram[20344] = 240;
// bram[20345] = 232;
// bram[20346] = 222;
// bram[20347] = 210;
// bram[20348] = 197;
// bram[20349] = 183;
// bram[20350] = 168;
// bram[20351] = 152;
// bram[20352] = 136;
// bram[20353] = 120;
// bram[20354] = 103;
// bram[20355] = 87;
// bram[20356] = 72;
// bram[20357] = 58;
// bram[20358] = 45;
// bram[20359] = 33;
// bram[20360] = 23;
// bram[20361] = 14;
// bram[20362] = 7;
// bram[20363] = 3;
// bram[20364] = 0;
// bram[20365] = 0;
// bram[20366] = 1;
// bram[20367] = 5;
// bram[20368] = 11;
// bram[20369] = 18;
// bram[20370] = 28;
// bram[20371] = 39;
// bram[20372] = 51;
// bram[20373] = 65;
// bram[20374] = 80;
// bram[20375] = 96;
// bram[20376] = 112;
// bram[20377] = 128;
// bram[20378] = 144;
// bram[20379] = 161;
// bram[20380] = 176;
// bram[20381] = 191;
// bram[20382] = 204;
// bram[20383] = 217;
// bram[20384] = 227;
// bram[20385] = 236;
// bram[20386] = 244;
// bram[20387] = 249;
// bram[20388] = 252;
// bram[20389] = 253;
// bram[20390] = 253;
// bram[20391] = 250;
// bram[20392] = 244;
// bram[20393] = 237;
// bram[20394] = 228;
// bram[20395] = 218;
// bram[20396] = 206;
// bram[20397] = 192;
// bram[20398] = 178;
// bram[20399] = 162;
// bram[20400] = 146;
// bram[20401] = 130;
// bram[20402] = 114;
// bram[20403] = 97;
// bram[20404] = 82;
// bram[20405] = 67;
// bram[20406] = 53;
// bram[20407] = 40;
// bram[20408] = 29;
// bram[20409] = 19;
// bram[20410] = 11;
// bram[20411] = 5;
// bram[20412] = 1;
// bram[20413] = 0;
// bram[20414] = 0;
// bram[20415] = 2;
// bram[20416] = 7;
// bram[20417] = 13;
// bram[20418] = 22;
// bram[20419] = 32;
// bram[20420] = 43;
// bram[20421] = 56;
// bram[20422] = 71;
// bram[20423] = 86;
// bram[20424] = 102;
// bram[20425] = 118;
// bram[20426] = 134;
// bram[20427] = 150;
// bram[20428] = 166;
// bram[20429] = 182;
// bram[20430] = 196;
// bram[20431] = 209;
// bram[20432] = 221;
// bram[20433] = 231;
// bram[20434] = 239;
// bram[20435] = 246;
// bram[20436] = 250;
// bram[20437] = 253;
// bram[20438] = 253;
// bram[20439] = 252;
// bram[20440] = 248;
// bram[20441] = 242;
// bram[20442] = 234;
// bram[20443] = 225;
// bram[20444] = 214;
// bram[20445] = 201;
// bram[20446] = 187;
// bram[20447] = 172;
// bram[20448] = 157;
// bram[20449] = 140;
// bram[20450] = 124;
// bram[20451] = 108;
// bram[20452] = 92;
// bram[20453] = 76;
// bram[20454] = 62;
// bram[20455] = 48;
// bram[20456] = 36;
// bram[20457] = 25;
// bram[20458] = 16;
// bram[20459] = 9;
// bram[20460] = 4;
// bram[20461] = 1;
// bram[20462] = 0;
// bram[20463] = 1;
// bram[20464] = 4;
// bram[20465] = 9;
// bram[20466] = 16;
// bram[20467] = 25;
// bram[20468] = 36;
// bram[20469] = 48;
// bram[20470] = 61;
// bram[20471] = 76;
// bram[20472] = 91;
// bram[20473] = 107;
// bram[20474] = 124;
// bram[20475] = 140;
// bram[20476] = 156;
// bram[20477] = 172;
// bram[20478] = 187;
// bram[20479] = 201;
// bram[20480] = 213;
// bram[20481] = 225;
// bram[20482] = 234;
// bram[20483] = 242;
// bram[20484] = 248;
// bram[20485] = 252;
// bram[20486] = 253;
// bram[20487] = 253;
// bram[20488] = 251;
// bram[20489] = 246;
// bram[20490] = 239;
// bram[20491] = 231;
// bram[20492] = 221;
// bram[20493] = 209;
// bram[20494] = 196;
// bram[20495] = 182;
// bram[20496] = 167;
// bram[20497] = 151;
// bram[20498] = 134;
// bram[20499] = 118;
// bram[20500] = 102;
// bram[20501] = 86;
// bram[20502] = 71;
// bram[20503] = 56;
// bram[20504] = 43;
// bram[20505] = 32;
// bram[20506] = 22;
// bram[20507] = 13;
// bram[20508] = 7;
// bram[20509] = 2;
// bram[20510] = 0;
// bram[20511] = 0;
// bram[20512] = 1;
// bram[20513] = 5;
// bram[20514] = 11;
// bram[20515] = 19;
// bram[20516] = 29;
// bram[20517] = 40;
// bram[20518] = 53;
// bram[20519] = 67;
// bram[20520] = 82;
// bram[20521] = 97;
// bram[20522] = 113;
// bram[20523] = 130;
// bram[20524] = 146;
// bram[20525] = 162;
// bram[20526] = 178;
// bram[20527] = 192;
// bram[20528] = 206;
// bram[20529] = 218;
// bram[20530] = 228;
// bram[20531] = 237;
// bram[20532] = 244;
// bram[20533] = 249;
// bram[20534] = 253;
// bram[20535] = 253;
// bram[20536] = 252;
// bram[20537] = 249;
// bram[20538] = 244;
// bram[20539] = 237;
// bram[20540] = 227;
// bram[20541] = 217;
// bram[20542] = 204;
// bram[20543] = 191;
// bram[20544] = 176;
// bram[20545] = 161;
// bram[20546] = 145;
// bram[20547] = 128;
// bram[20548] = 112;
// bram[20549] = 96;
// bram[20550] = 80;
// bram[20551] = 65;
// bram[20552] = 52;
// bram[20553] = 39;
// bram[20554] = 28;
// bram[20555] = 18;
// bram[20556] = 11;
// bram[20557] = 5;
// bram[20558] = 1;
// bram[20559] = 0;
// bram[20560] = 0;
// bram[20561] = 3;
// bram[20562] = 7;
// bram[20563] = 14;
// bram[20564] = 22;
// bram[20565] = 33;
// bram[20566] = 45;
// bram[20567] = 58;
// bram[20568] = 72;
// bram[20569] = 87;
// bram[20570] = 103;
// bram[20571] = 119;
// bram[20572] = 136;
// bram[20573] = 152;
// bram[20574] = 168;
// bram[20575] = 183;
// bram[20576] = 197;
// bram[20577] = 210;
// bram[20578] = 222;
// bram[20579] = 232;
// bram[20580] = 240;
// bram[20581] = 246;
// bram[20582] = 251;
// bram[20583] = 253;
// bram[20584] = 253;
// bram[20585] = 251;
// bram[20586] = 247;
// bram[20587] = 241;
// bram[20588] = 233;
// bram[20589] = 224;
// bram[20590] = 212;
// bram[20591] = 200;
// bram[20592] = 186;
// bram[20593] = 171;
// bram[20594] = 155;
// bram[20595] = 139;
// bram[20596] = 122;
// bram[20597] = 106;
// bram[20598] = 90;
// bram[20599] = 75;
// bram[20600] = 60;
// bram[20601] = 47;
// bram[20602] = 35;
// bram[20603] = 24;
// bram[20604] = 15;
// bram[20605] = 8;
// bram[20606] = 3;
// bram[20607] = 0;
// bram[20608] = 0;
// bram[20609] = 1;
// bram[20610] = 4;
// bram[20611] = 10;
// bram[20612] = 17;
// bram[20613] = 26;
// bram[20614] = 37;
// bram[20615] = 49;
// bram[20616] = 63;
// bram[20617] = 78;
// bram[20618] = 93;
// bram[20619] = 109;
// bram[20620] = 126;
// bram[20621] = 142;
// bram[20622] = 158;
// bram[20623] = 174;
// bram[20624] = 188;
// bram[20625] = 202;
// bram[20626] = 215;
// bram[20627] = 226;
// bram[20628] = 235;
// bram[20629] = 243;
// bram[20630] = 248;
// bram[20631] = 252;
// bram[20632] = 253;
// bram[20633] = 253;
// bram[20634] = 250;
// bram[20635] = 245;
// bram[20636] = 239;
// bram[20637] = 230;
// bram[20638] = 220;
// bram[20639] = 208;
// bram[20640] = 195;
// bram[20641] = 180;
// bram[20642] = 165;
// bram[20643] = 149;
// bram[20644] = 133;
// bram[20645] = 116;
// bram[20646] = 100;
// bram[20647] = 84;
// bram[20648] = 69;
// bram[20649] = 55;
// bram[20650] = 42;
// bram[20651] = 31;
// bram[20652] = 21;
// bram[20653] = 13;
// bram[20654] = 6;
// bram[20655] = 2;
// bram[20656] = 0;
// bram[20657] = 0;
// bram[20658] = 2;
// bram[20659] = 6;
// bram[20660] = 12;
// bram[20661] = 20;
// bram[20662] = 30;
// bram[20663] = 41;
// bram[20664] = 54;
// bram[20665] = 68;
// bram[20666] = 83;
// bram[20667] = 99;
// bram[20668] = 115;
// bram[20669] = 132;
// bram[20670] = 148;
// bram[20671] = 164;
// bram[20672] = 179;
// bram[20673] = 194;
// bram[20674] = 207;
// bram[20675] = 219;
// bram[20676] = 229;
// bram[20677] = 238;
// bram[20678] = 245;
// bram[20679] = 250;
// bram[20680] = 253;
// bram[20681] = 253;
// bram[20682] = 252;
// bram[20683] = 249;
// bram[20684] = 243;
// bram[20685] = 236;
// bram[20686] = 226;
// bram[20687] = 215;
// bram[20688] = 203;
// bram[20689] = 189;
// bram[20690] = 175;
// bram[20691] = 159;
// bram[20692] = 143;
// bram[20693] = 127;
// bram[20694] = 110;
// bram[20695] = 94;
// bram[20696] = 79;
// bram[20697] = 64;
// bram[20698] = 50;
// bram[20699] = 38;
// bram[20700] = 27;
// bram[20701] = 17;
// bram[20702] = 10;
// bram[20703] = 4;
// bram[20704] = 1;
// bram[20705] = 0;
// bram[20706] = 0;
// bram[20707] = 3;
// bram[20708] = 8;
// bram[20709] = 15;
// bram[20710] = 23;
// bram[20711] = 34;
// bram[20712] = 46;
// bram[20713] = 59;
// bram[20714] = 74;
// bram[20715] = 89;
// bram[20716] = 105;
// bram[20717] = 121;
// bram[20718] = 138;
// bram[20719] = 154;
// bram[20720] = 170;
// bram[20721] = 185;
// bram[20722] = 199;
// bram[20723] = 211;
// bram[20724] = 223;
// bram[20725] = 233;
// bram[20726] = 241;
// bram[20727] = 247;
// bram[20728] = 251;
// bram[20729] = 253;
// bram[20730] = 253;
// bram[20731] = 251;
// bram[20732] = 247;
// bram[20733] = 241;
// bram[20734] = 232;
// bram[20735] = 223;
// bram[20736] = 211;
// bram[20737] = 198;
// bram[20738] = 184;
// bram[20739] = 169;
// bram[20740] = 153;
// bram[20741] = 137;
// bram[20742] = 121;
// bram[20743] = 104;
// bram[20744] = 88;
// bram[20745] = 73;
// bram[20746] = 59;
// bram[20747] = 45;
// bram[20748] = 34;
// bram[20749] = 23;
// bram[20750] = 14;
// bram[20751] = 8;
// bram[20752] = 3;
// bram[20753] = 0;
// bram[20754] = 0;
// bram[20755] = 1;
// bram[20756] = 5;
// bram[20757] = 10;
// bram[20758] = 18;
// bram[20759] = 27;
// bram[20760] = 38;
// bram[20761] = 51;
// bram[20762] = 64;
// bram[20763] = 79;
// bram[20764] = 95;
// bram[20765] = 111;
// bram[20766] = 127;
// bram[20767] = 144;
// bram[20768] = 160;
// bram[20769] = 175;
// bram[20770] = 190;
// bram[20771] = 204;
// bram[20772] = 216;
// bram[20773] = 227;
// bram[20774] = 236;
// bram[20775] = 243;
// bram[20776] = 249;
// bram[20777] = 252;
// bram[20778] = 253;
// bram[20779] = 253;
// bram[20780] = 250;
// bram[20781] = 245;
// bram[20782] = 238;
// bram[20783] = 229;
// bram[20784] = 219;
// bram[20785] = 206;
// bram[20786] = 193;
// bram[20787] = 179;
// bram[20788] = 163;
// bram[20789] = 147;
// bram[20790] = 131;
// bram[20791] = 115;
// bram[20792] = 98;
// bram[20793] = 83;
// bram[20794] = 68;
// bram[20795] = 54;
// bram[20796] = 41;
// bram[20797] = 30;
// bram[20798] = 20;
// bram[20799] = 12;
// bram[20800] = 6;
// bram[20801] = 2;
// bram[20802] = 0;
// bram[20803] = 0;
// bram[20804] = 2;
// bram[20805] = 6;
// bram[20806] = 13;
// bram[20807] = 21;
// bram[20808] = 31;
// bram[20809] = 43;
// bram[20810] = 56;
// bram[20811] = 70;
// bram[20812] = 85;
// bram[20813] = 101;
// bram[20814] = 117;
// bram[20815] = 133;
// bram[20816] = 150;
// bram[20817] = 165;
// bram[20818] = 181;
// bram[20819] = 195;
// bram[20820] = 208;
// bram[20821] = 220;
// bram[20822] = 230;
// bram[20823] = 239;
// bram[20824] = 246;
// bram[20825] = 250;
// bram[20826] = 253;
// bram[20827] = 253;
// bram[20828] = 252;
// bram[20829] = 248;
// bram[20830] = 242;
// bram[20831] = 235;
// bram[20832] = 225;
// bram[20833] = 214;
// bram[20834] = 202;
// bram[20835] = 188;
// bram[20836] = 173;
// bram[20837] = 157;
// bram[20838] = 141;
// bram[20839] = 125;
// bram[20840] = 109;
// bram[20841] = 93;
// bram[20842] = 77;
// bram[20843] = 62;
// bram[20844] = 49;
// bram[20845] = 37;
// bram[20846] = 26;
// bram[20847] = 17;
// bram[20848] = 9;
// bram[20849] = 4;
// bram[20850] = 1;
// bram[20851] = 0;
// bram[20852] = 0;
// bram[20853] = 3;
// bram[20854] = 9;
// bram[20855] = 16;
// bram[20856] = 24;
// bram[20857] = 35;
// bram[20858] = 47;
// bram[20859] = 61;
// bram[20860] = 75;
// bram[20861] = 91;
// bram[20862] = 107;
// bram[20863] = 123;
// bram[20864] = 139;
// bram[20865] = 155;
// bram[20866] = 171;
// bram[20867] = 186;
// bram[20868] = 200;
// bram[20869] = 213;
// bram[20870] = 224;
// bram[20871] = 234;
// bram[20872] = 242;
// bram[20873] = 248;
// bram[20874] = 251;
// bram[20875] = 253;
// bram[20876] = 253;
// bram[20877] = 251;
// bram[20878] = 246;
// bram[20879] = 240;
// bram[20880] = 232;
// bram[20881] = 221;
// bram[20882] = 210;
// bram[20883] = 197;
// bram[20884] = 183;
// bram[20885] = 167;
// bram[20886] = 152;
// bram[20887] = 135;
// bram[20888] = 119;
// bram[20889] = 103;
// bram[20890] = 87;
// bram[20891] = 72;
// bram[20892] = 57;
// bram[20893] = 44;
// bram[20894] = 32;
// bram[20895] = 22;
// bram[20896] = 14;
// bram[20897] = 7;
// bram[20898] = 3;
// bram[20899] = 0;
// bram[20900] = 0;
// bram[20901] = 1;
// bram[20902] = 5;
// bram[20903] = 11;
// bram[20904] = 19;
// bram[20905] = 28;
// bram[20906] = 39;
// bram[20907] = 52;
// bram[20908] = 66;
// bram[20909] = 81;
// bram[20910] = 96;
// bram[20911] = 113;
// bram[20912] = 129;
// bram[20913] = 145;
// bram[20914] = 161;
// bram[20915] = 177;
// bram[20916] = 191;
// bram[20917] = 205;
// bram[20918] = 217;
// bram[20919] = 228;
// bram[20920] = 237;
// bram[20921] = 244;
// bram[20922] = 249;
// bram[20923] = 252;
// bram[20924] = 253;
// bram[20925] = 252;
// bram[20926] = 249;
// bram[20927] = 244;
// bram[20928] = 237;
// bram[20929] = 228;
// bram[20930] = 217;
// bram[20931] = 205;
// bram[20932] = 192;
// bram[20933] = 177;
// bram[20934] = 162;
// bram[20935] = 146;
// bram[20936] = 129;
// bram[20937] = 113;
// bram[20938] = 97;
// bram[20939] = 81;
// bram[20940] = 66;
// bram[20941] = 52;
// bram[20942] = 40;
// bram[20943] = 28;
// bram[20944] = 19;
// bram[20945] = 11;
// bram[20946] = 5;
// bram[20947] = 1;
// bram[20948] = 0;
// bram[20949] = 0;
// bram[20950] = 2;
// bram[20951] = 7;
// bram[20952] = 14;
// bram[20953] = 22;
// bram[20954] = 32;
// bram[20955] = 44;
// bram[20956] = 57;
// bram[20957] = 71;
// bram[20958] = 86;
// bram[20959] = 102;
// bram[20960] = 119;
// bram[20961] = 135;
// bram[20962] = 151;
// bram[20963] = 167;
// bram[20964] = 182;
// bram[20965] = 196;
// bram[20966] = 210;
// bram[20967] = 221;
// bram[20968] = 231;
// bram[20969] = 240;
// bram[20970] = 246;
// bram[20971] = 251;
// bram[20972] = 253;
// bram[20973] = 253;
// bram[20974] = 252;
// bram[20975] = 248;
// bram[20976] = 242;
// bram[20977] = 234;
// bram[20978] = 224;
// bram[20979] = 213;
// bram[20980] = 200;
// bram[20981] = 186;
// bram[20982] = 171;
// bram[20983] = 156;
// bram[20984] = 140;
// bram[20985] = 123;
// bram[20986] = 107;
// bram[20987] = 91;
// bram[20988] = 76;
// bram[20989] = 61;
// bram[20990] = 47;
// bram[20991] = 35;
// bram[20992] = 25;
// bram[20993] = 16;
// bram[20994] = 9;
// bram[20995] = 4;
// bram[20996] = 0;
// bram[20997] = 0;
// bram[20998] = 1;
// bram[20999] = 4;
// bram[21000] = 9;
// bram[21001] = 16;
// bram[21002] = 25;
// bram[21003] = 36;
// bram[21004] = 49;
// bram[21005] = 62;
// bram[21006] = 77;
// bram[21007] = 92;
// bram[21008] = 108;
// bram[21009] = 125;
// bram[21010] = 141;
// bram[21011] = 157;
// bram[21012] = 173;
// bram[21013] = 188;
// bram[21014] = 201;
// bram[21015] = 214;
// bram[21016] = 225;
// bram[21017] = 235;
// bram[21018] = 242;
// bram[21019] = 248;
// bram[21020] = 252;
// bram[21021] = 253;
// bram[21022] = 253;
// bram[21023] = 250;
// bram[21024] = 246;
// bram[21025] = 239;
// bram[21026] = 231;
// bram[21027] = 220;
// bram[21028] = 209;
// bram[21029] = 195;
// bram[21030] = 181;
// bram[21031] = 166;
// bram[21032] = 150;
// bram[21033] = 134;
// bram[21034] = 117;
// bram[21035] = 101;
// bram[21036] = 85;
// bram[21037] = 70;
// bram[21038] = 56;
// bram[21039] = 43;
// bram[21040] = 31;
// bram[21041] = 21;
// bram[21042] = 13;
// bram[21043] = 7;
// bram[21044] = 2;
// bram[21045] = 0;
// bram[21046] = 0;
// bram[21047] = 2;
// bram[21048] = 6;
// bram[21049] = 12;
// bram[21050] = 20;
// bram[21051] = 29;
// bram[21052] = 41;
// bram[21053] = 53;
// bram[21054] = 67;
// bram[21055] = 82;
// bram[21056] = 98;
// bram[21057] = 114;
// bram[21058] = 131;
// bram[21059] = 147;
// bram[21060] = 163;
// bram[21061] = 178;
// bram[21062] = 193;
// bram[21063] = 206;
// bram[21064] = 218;
// bram[21065] = 229;
// bram[21066] = 238;
// bram[21067] = 245;
// bram[21068] = 250;
// bram[21069] = 253;
// bram[21070] = 253;
// bram[21071] = 252;
// bram[21072] = 249;
// bram[21073] = 244;
// bram[21074] = 236;
// bram[21075] = 227;
// bram[21076] = 216;
// bram[21077] = 204;
// bram[21078] = 190;
// bram[21079] = 176;
// bram[21080] = 160;
// bram[21081] = 144;
// bram[21082] = 128;
// bram[21083] = 111;
// bram[21084] = 95;
// bram[21085] = 80;
// bram[21086] = 65;
// bram[21087] = 51;
// bram[21088] = 38;
// bram[21089] = 27;
// bram[21090] = 18;
// bram[21091] = 10;
// bram[21092] = 5;
// bram[21093] = 1;
// bram[21094] = 0;
// bram[21095] = 0;
// bram[21096] = 3;
// bram[21097] = 8;
// bram[21098] = 14;
// bram[21099] = 23;
// bram[21100] = 33;
// bram[21101] = 45;
// bram[21102] = 58;
// bram[21103] = 73;
// bram[21104] = 88;
// bram[21105] = 104;
// bram[21106] = 120;
// bram[21107] = 137;
// bram[21108] = 153;
// bram[21109] = 169;
// bram[21110] = 184;
// bram[21111] = 198;
// bram[21112] = 211;
// bram[21113] = 222;
// bram[21114] = 232;
// bram[21115] = 240;
// bram[21116] = 247;
// bram[21117] = 251;
// bram[21118] = 253;
// bram[21119] = 253;
// bram[21120] = 251;
// bram[21121] = 247;
// bram[21122] = 241;
// bram[21123] = 233;
// bram[21124] = 223;
// bram[21125] = 212;
// bram[21126] = 199;
// bram[21127] = 185;
// bram[21128] = 170;
// bram[21129] = 154;
// bram[21130] = 138;
// bram[21131] = 122;
// bram[21132] = 105;
// bram[21133] = 89;
// bram[21134] = 74;
// bram[21135] = 60;
// bram[21136] = 46;
// bram[21137] = 34;
// bram[21138] = 24;
// bram[21139] = 15;
// bram[21140] = 8;
// bram[21141] = 3;
// bram[21142] = 0;
// bram[21143] = 0;
// bram[21144] = 1;
// bram[21145] = 4;
// bram[21146] = 10;
// bram[21147] = 17;
// bram[21148] = 27;
// bram[21149] = 37;
// bram[21150] = 50;
// bram[21151] = 64;
// bram[21152] = 78;
// bram[21153] = 94;
// bram[21154] = 110;
// bram[21155] = 126;
// bram[21156] = 143;
// bram[21157] = 159;
// bram[21158] = 174;
// bram[21159] = 189;
// bram[21160] = 203;
// bram[21161] = 215;
// bram[21162] = 226;
// bram[21163] = 235;
// bram[21164] = 243;
// bram[21165] = 249;
// bram[21166] = 252;
// bram[21167] = 253;
// bram[21168] = 253;
// bram[21169] = 250;
// bram[21170] = 245;
// bram[21171] = 238;
// bram[21172] = 230;
// bram[21173] = 219;
// bram[21174] = 207;
// bram[21175] = 194;
// bram[21176] = 179;
// bram[21177] = 164;
// bram[21178] = 148;
// bram[21179] = 132;
// bram[21180] = 116;
// bram[21181] = 99;
// bram[21182] = 84;
// bram[21183] = 69;
// bram[21184] = 54;
// bram[21185] = 42;
// bram[21186] = 30;
// bram[21187] = 20;
// bram[21188] = 12;
// bram[21189] = 6;
// bram[21190] = 2;
// bram[21191] = 0;
// bram[21192] = 0;
// bram[21193] = 2;
// bram[21194] = 6;
// bram[21195] = 12;
// bram[21196] = 20;
// bram[21197] = 30;
// bram[21198] = 42;
// bram[21199] = 55;
// bram[21200] = 69;
// bram[21201] = 84;
// bram[21202] = 100;
// bram[21203] = 116;
// bram[21204] = 132;
// bram[21205] = 149;
// bram[21206] = 165;
// bram[21207] = 180;
// bram[21208] = 194;
// bram[21209] = 207;
// bram[21210] = 219;
// bram[21211] = 230;
// bram[21212] = 238;
// bram[21213] = 245;
// bram[21214] = 250;
// bram[21215] = 253;
// bram[21216] = 253;
// bram[21217] = 252;
// bram[21218] = 248;
// bram[21219] = 243;
// bram[21220] = 235;
// bram[21221] = 226;
// bram[21222] = 215;
// bram[21223] = 202;
// bram[21224] = 189;
// bram[21225] = 174;
// bram[21226] = 158;
// bram[21227] = 142;
// bram[21228] = 126;
// bram[21229] = 110;
// bram[21230] = 93;
// bram[21231] = 78;
// bram[21232] = 63;
// bram[21233] = 50;
// bram[21234] = 37;
// bram[21235] = 26;
// bram[21236] = 17;
// bram[21237] = 10;
// bram[21238] = 4;
// bram[21239] = 1;
// bram[21240] = 0;
// bram[21241] = 0;
// bram[21242] = 3;
// bram[21243] = 8;
// bram[21244] = 15;
// bram[21245] = 24;
// bram[21246] = 34;
// bram[21247] = 46;
// bram[21248] = 60;
// bram[21249] = 74;
// bram[21250] = 90;
// bram[21251] = 106;
// bram[21252] = 122;
// bram[21253] = 138;
// bram[21254] = 154;
// bram[21255] = 170;
// bram[21256] = 185;
// bram[21257] = 199;
// bram[21258] = 212;
// bram[21259] = 223;
// bram[21260] = 233;
// bram[21261] = 241;
// bram[21262] = 247;
// bram[21263] = 251;
// bram[21264] = 253;
// bram[21265] = 253;
// bram[21266] = 251;
// bram[21267] = 247;
// bram[21268] = 240;
// bram[21269] = 232;
// bram[21270] = 222;
// bram[21271] = 211;
// bram[21272] = 198;
// bram[21273] = 183;
// bram[21274] = 168;
// bram[21275] = 152;
// bram[21276] = 136;
// bram[21277] = 120;
// bram[21278] = 104;
// bram[21279] = 88;
// bram[21280] = 72;
// bram[21281] = 58;
// bram[21282] = 45;
// bram[21283] = 33;
// bram[21284] = 23;
// bram[21285] = 14;
// bram[21286] = 7;
// bram[21287] = 3;
// bram[21288] = 0;
// bram[21289] = 0;
// bram[21290] = 1;
// bram[21291] = 5;
// bram[21292] = 11;
// bram[21293] = 18;
// bram[21294] = 28;
// bram[21295] = 39;
// bram[21296] = 51;
// bram[21297] = 65;
// bram[21298] = 80;
// bram[21299] = 95;
// bram[21300] = 112;
// bram[21301] = 128;
// bram[21302] = 144;
// bram[21303] = 160;
// bram[21304] = 176;
// bram[21305] = 191;
// bram[21306] = 204;
// bram[21307] = 216;
// bram[21308] = 227;
// bram[21309] = 236;
// bram[21310] = 244;
// bram[21311] = 249;
// bram[21312] = 252;
// bram[21313] = 253;
// bram[21314] = 253;
// bram[21315] = 250;
// bram[21316] = 245;
// bram[21317] = 237;
// bram[21318] = 229;
// bram[21319] = 218;
// bram[21320] = 206;
// bram[21321] = 192;
// bram[21322] = 178;
// bram[21323] = 163;
// bram[21324] = 147;
// bram[21325] = 130;
// bram[21326] = 114;
// bram[21327] = 98;
// bram[21328] = 82;
// bram[21329] = 67;
// bram[21330] = 53;
// bram[21331] = 40;
// bram[21332] = 29;
// bram[21333] = 19;
// bram[21334] = 11;
// bram[21335] = 5;
// bram[21336] = 2;
// bram[21337] = 0;
// bram[21338] = 0;
// bram[21339] = 2;
// bram[21340] = 7;
// bram[21341] = 13;
// bram[21342] = 21;
// bram[21343] = 31;
// bram[21344] = 43;
// bram[21345] = 56;
// bram[21346] = 70;
// bram[21347] = 86;
// bram[21348] = 101;
// bram[21349] = 118;
// bram[21350] = 134;
// bram[21351] = 150;
// bram[21352] = 166;
// bram[21353] = 181;
// bram[21354] = 196;
// bram[21355] = 209;
// bram[21356] = 221;
// bram[21357] = 231;
// bram[21358] = 239;
// bram[21359] = 246;
// bram[21360] = 250;
// bram[21361] = 253;
// bram[21362] = 253;
// bram[21363] = 252;
// bram[21364] = 248;
// bram[21365] = 242;
// bram[21366] = 234;
// bram[21367] = 225;
// bram[21368] = 214;
// bram[21369] = 201;
// bram[21370] = 187;
// bram[21371] = 172;
// bram[21372] = 157;
// bram[21373] = 141;
// bram[21374] = 124;
// bram[21375] = 108;
// bram[21376] = 92;
// bram[21377] = 76;
// bram[21378] = 62;
// bram[21379] = 48;
// bram[21380] = 36;
// bram[21381] = 25;
// bram[21382] = 16;
// bram[21383] = 9;
// bram[21384] = 4;
// bram[21385] = 1;
// bram[21386] = 0;
// bram[21387] = 1;
// bram[21388] = 4;
// bram[21389] = 9;
// bram[21390] = 16;
// bram[21391] = 25;
// bram[21392] = 36;
// bram[21393] = 48;
// bram[21394] = 61;
// bram[21395] = 76;
// bram[21396] = 91;
// bram[21397] = 107;
// bram[21398] = 124;
// bram[21399] = 140;
// bram[21400] = 156;
// bram[21401] = 172;
// bram[21402] = 187;
// bram[21403] = 201;
// bram[21404] = 213;
// bram[21405] = 225;
// bram[21406] = 234;
// bram[21407] = 242;
// bram[21408] = 248;
// bram[21409] = 252;
// bram[21410] = 253;
// bram[21411] = 253;
// bram[21412] = 251;
// bram[21413] = 246;
// bram[21414] = 240;
// bram[21415] = 231;
// bram[21416] = 221;
// bram[21417] = 209;
// bram[21418] = 196;
// bram[21419] = 182;
// bram[21420] = 167;
// bram[21421] = 151;
// bram[21422] = 135;
// bram[21423] = 118;
// bram[21424] = 102;
// bram[21425] = 86;
// bram[21426] = 71;
// bram[21427] = 57;
// bram[21428] = 44;
// bram[21429] = 32;
// bram[21430] = 22;
// bram[21431] = 13;
// bram[21432] = 7;
// bram[21433] = 2;
// bram[21434] = 0;
// bram[21435] = 0;
// bram[21436] = 1;
// bram[21437] = 5;
// bram[21438] = 11;
// bram[21439] = 19;
// bram[21440] = 29;
// bram[21441] = 40;
// bram[21442] = 53;
// bram[21443] = 67;
// bram[21444] = 81;
// bram[21445] = 97;
// bram[21446] = 113;
// bram[21447] = 130;
// bram[21448] = 146;
// bram[21449] = 162;
// bram[21450] = 177;
// bram[21451] = 192;
// bram[21452] = 205;
// bram[21453] = 218;
// bram[21454] = 228;
// bram[21455] = 237;
// bram[21456] = 244;
// bram[21457] = 249;
// bram[21458] = 253;
// bram[21459] = 253;
// bram[21460] = 252;
// bram[21461] = 249;
// bram[21462] = 244;
// bram[21463] = 237;
// bram[21464] = 228;
// bram[21465] = 217;
// bram[21466] = 205;
// bram[21467] = 191;
// bram[21468] = 176;
// bram[21469] = 161;
// bram[21470] = 145;
// bram[21471] = 129;
// bram[21472] = 112;
// bram[21473] = 96;
// bram[21474] = 80;
// bram[21475] = 66;
// bram[21476] = 52;
// bram[21477] = 39;
// bram[21478] = 28;
// bram[21479] = 18;
// bram[21480] = 11;
// bram[21481] = 5;
// bram[21482] = 1;
// bram[21483] = 0;
// bram[21484] = 0;
// bram[21485] = 3;
// bram[21486] = 7;
// bram[21487] = 14;
// bram[21488] = 22;
// bram[21489] = 33;
// bram[21490] = 44;
// bram[21491] = 58;
// bram[21492] = 72;
// bram[21493] = 87;
// bram[21494] = 103;
// bram[21495] = 119;
// bram[21496] = 136;
// bram[21497] = 152;
// bram[21498] = 168;
// bram[21499] = 183;
// bram[21500] = 197;
// bram[21501] = 210;
// bram[21502] = 222;
// bram[21503] = 232;
// bram[21504] = 240;
// bram[21505] = 246;
// bram[21506] = 251;
// bram[21507] = 253;
// bram[21508] = 253;
// bram[21509] = 251;
// bram[21510] = 247;
// bram[21511] = 241;
// bram[21512] = 234;
// bram[21513] = 224;
// bram[21514] = 212;
// bram[21515] = 200;
// bram[21516] = 186;
// bram[21517] = 171;
// bram[21518] = 155;
// bram[21519] = 139;
// bram[21520] = 123;
// bram[21521] = 106;
// bram[21522] = 90;
// bram[21523] = 75;
// bram[21524] = 60;
// bram[21525] = 47;
// bram[21526] = 35;
// bram[21527] = 24;
// bram[21528] = 15;
// bram[21529] = 8;
// bram[21530] = 3;
// bram[21531] = 0;
// bram[21532] = 0;
// bram[21533] = 1;
// bram[21534] = 4;
// bram[21535] = 9;
// bram[21536] = 17;
// bram[21537] = 26;
// bram[21538] = 37;
// bram[21539] = 49;
// bram[21540] = 63;
// bram[21541] = 77;
// bram[21542] = 93;
// bram[21543] = 109;
// bram[21544] = 125;
// bram[21545] = 142;
// bram[21546] = 158;
// bram[21547] = 173;
// bram[21548] = 188;
// bram[21549] = 202;
// bram[21550] = 215;
// bram[21551] = 226;
// bram[21552] = 235;
// bram[21553] = 243;
// bram[21554] = 248;
// bram[21555] = 252;
// bram[21556] = 253;
// bram[21557] = 253;
// bram[21558] = 250;
// bram[21559] = 245;
// bram[21560] = 239;
// bram[21561] = 230;
// bram[21562] = 220;
// bram[21563] = 208;
// bram[21564] = 195;
// bram[21565] = 180;
// bram[21566] = 165;
// bram[21567] = 149;
// bram[21568] = 133;
// bram[21569] = 116;
// bram[21570] = 100;
// bram[21571] = 84;
// bram[21572] = 69;
// bram[21573] = 55;
// bram[21574] = 42;
// bram[21575] = 31;
// bram[21576] = 21;
// bram[21577] = 13;
// bram[21578] = 6;
// bram[21579] = 2;
// bram[21580] = 0;
// bram[21581] = 0;
// bram[21582] = 2;
// bram[21583] = 6;
// bram[21584] = 12;
// bram[21585] = 20;
// bram[21586] = 30;
// bram[21587] = 41;
// bram[21588] = 54;
// bram[21589] = 68;
// bram[21590] = 83;
// bram[21591] = 99;
// bram[21592] = 115;
// bram[21593] = 131;
// bram[21594] = 148;
// bram[21595] = 164;
// bram[21596] = 179;
// bram[21597] = 193;
// bram[21598] = 207;
// bram[21599] = 219;
// bram[21600] = 229;
// bram[21601] = 238;
// bram[21602] = 245;
// bram[21603] = 250;
// bram[21604] = 253;
// bram[21605] = 253;
// bram[21606] = 252;
// bram[21607] = 249;
// bram[21608] = 243;
// bram[21609] = 236;
// bram[21610] = 227;
// bram[21611] = 216;
// bram[21612] = 203;
// bram[21613] = 190;
// bram[21614] = 175;
// bram[21615] = 159;
// bram[21616] = 143;
// bram[21617] = 127;
// bram[21618] = 110;
// bram[21619] = 94;
// bram[21620] = 79;
// bram[21621] = 64;
// bram[21622] = 50;
// bram[21623] = 38;
// bram[21624] = 27;
// bram[21625] = 18;
// bram[21626] = 10;
// bram[21627] = 5;
// bram[21628] = 1;
// bram[21629] = 0;
// bram[21630] = 0;
// bram[21631] = 3;
// bram[21632] = 8;
// bram[21633] = 15;
// bram[21634] = 23;
// bram[21635] = 34;
// bram[21636] = 46;
// bram[21637] = 59;
// bram[21638] = 73;
// bram[21639] = 89;
// bram[21640] = 105;
// bram[21641] = 121;
// bram[21642] = 137;
// bram[21643] = 154;
// bram[21644] = 169;
// bram[21645] = 184;
// bram[21646] = 198;
// bram[21647] = 211;
// bram[21648] = 223;
// bram[21649] = 233;
// bram[21650] = 241;
// bram[21651] = 247;
// bram[21652] = 251;
// bram[21653] = 253;
// bram[21654] = 253;
// bram[21655] = 251;
// bram[21656] = 247;
// bram[21657] = 241;
// bram[21658] = 233;
// bram[21659] = 223;
// bram[21660] = 211;
// bram[21661] = 198;
// bram[21662] = 184;
// bram[21663] = 169;
// bram[21664] = 153;
// bram[21665] = 137;
// bram[21666] = 121;
// bram[21667] = 105;
// bram[21668] = 89;
// bram[21669] = 73;
// bram[21670] = 59;
// bram[21671] = 46;
// bram[21672] = 34;
// bram[21673] = 23;
// bram[21674] = 15;
// bram[21675] = 8;
// bram[21676] = 3;
// bram[21677] = 0;
// bram[21678] = 0;
// bram[21679] = 1;
// bram[21680] = 5;
// bram[21681] = 10;
// bram[21682] = 18;
// bram[21683] = 27;
// bram[21684] = 38;
// bram[21685] = 50;
// bram[21686] = 64;
// bram[21687] = 79;
// bram[21688] = 95;
// bram[21689] = 111;
// bram[21690] = 127;
// bram[21691] = 143;
// bram[21692] = 159;
// bram[21693] = 175;
// bram[21694] = 190;
// bram[21695] = 203;
// bram[21696] = 216;
// bram[21697] = 227;
// bram[21698] = 236;
// bram[21699] = 243;
// bram[21700] = 249;
// bram[21701] = 252;
// bram[21702] = 253;
// bram[21703] = 253;
// bram[21704] = 250;
// bram[21705] = 245;
// bram[21706] = 238;
// bram[21707] = 229;
// bram[21708] = 219;
// bram[21709] = 207;
// bram[21710] = 193;
// bram[21711] = 179;
// bram[21712] = 163;
// bram[21713] = 147;
// bram[21714] = 131;
// bram[21715] = 115;
// bram[21716] = 99;
// bram[21717] = 83;
// bram[21718] = 68;
// bram[21719] = 54;
// bram[21720] = 41;
// bram[21721] = 30;
// bram[21722] = 20;
// bram[21723] = 12;
// bram[21724] = 6;
// bram[21725] = 2;
// bram[21726] = 0;
// bram[21727] = 0;
// bram[21728] = 2;
// bram[21729] = 6;
// bram[21730] = 13;
// bram[21731] = 21;
// bram[21732] = 31;
// bram[21733] = 42;
// bram[21734] = 55;
// bram[21735] = 70;
// bram[21736] = 85;
// bram[21737] = 100;
// bram[21738] = 117;
// bram[21739] = 133;
// bram[21740] = 149;
// bram[21741] = 165;
// bram[21742] = 180;
// bram[21743] = 195;
// bram[21744] = 208;
// bram[21745] = 220;
// bram[21746] = 230;
// bram[21747] = 239;
// bram[21748] = 246;
// bram[21749] = 250;
// bram[21750] = 253;
// bram[21751] = 253;
// bram[21752] = 252;
// bram[21753] = 248;
// bram[21754] = 243;
// bram[21755] = 235;
// bram[21756] = 225;
// bram[21757] = 214;
// bram[21758] = 202;
// bram[21759] = 188;
// bram[21760] = 173;
// bram[21761] = 158;
// bram[21762] = 142;
// bram[21763] = 125;
// bram[21764] = 109;
// bram[21765] = 93;
// bram[21766] = 77;
// bram[21767] = 63;
// bram[21768] = 49;
// bram[21769] = 37;
// bram[21770] = 26;
// bram[21771] = 17;
// bram[21772] = 9;
// bram[21773] = 4;
// bram[21774] = 1;
// bram[21775] = 0;
// bram[21776] = 0;
// bram[21777] = 3;
// bram[21778] = 8;
// bram[21779] = 15;
// bram[21780] = 24;
// bram[21781] = 35;
// bram[21782] = 47;
// bram[21783] = 60;
// bram[21784] = 75;
// bram[21785] = 90;
// bram[21786] = 106;
// bram[21787] = 123;
// bram[21788] = 139;
// bram[21789] = 155;
// bram[21790] = 171;
// bram[21791] = 186;
// bram[21792] = 200;
// bram[21793] = 213;
// bram[21794] = 224;
// bram[21795] = 234;
// bram[21796] = 241;
// bram[21797] = 247;
// bram[21798] = 251;
// bram[21799] = 253;
// bram[21800] = 253;
// bram[21801] = 251;
// bram[21802] = 246;
// bram[21803] = 240;
// bram[21804] = 232;
// bram[21805] = 222;
// bram[21806] = 210;
// bram[21807] = 197;
// bram[21808] = 183;
// bram[21809] = 168;
// bram[21810] = 152;
// bram[21811] = 136;
// bram[21812] = 119;
// bram[21813] = 103;
// bram[21814] = 87;
// bram[21815] = 72;
// bram[21816] = 57;
// bram[21817] = 44;
// bram[21818] = 32;
// bram[21819] = 22;
// bram[21820] = 14;
// bram[21821] = 7;
// bram[21822] = 3;
// bram[21823] = 0;
// bram[21824] = 0;
// bram[21825] = 1;
// bram[21826] = 5;
// bram[21827] = 11;
// bram[21828] = 19;
// bram[21829] = 28;
// bram[21830] = 39;
// bram[21831] = 52;
// bram[21832] = 66;
// bram[21833] = 81;
// bram[21834] = 96;
// bram[21835] = 112;
// bram[21836] = 129;
// bram[21837] = 145;
// bram[21838] = 161;
// bram[21839] = 177;
// bram[21840] = 191;
// bram[21841] = 205;
// bram[21842] = 217;
// bram[21843] = 228;
// bram[21844] = 237;
// bram[21845] = 244;
// bram[21846] = 249;
// bram[21847] = 252;
// bram[21848] = 253;
// bram[21849] = 252;
// bram[21850] = 249;
// bram[21851] = 244;
// bram[21852] = 237;
// bram[21853] = 228;
// bram[21854] = 217;
// bram[21855] = 205;
// bram[21856] = 192;
// bram[21857] = 177;
// bram[21858] = 162;
// bram[21859] = 146;
// bram[21860] = 129;
// bram[21861] = 113;
// bram[21862] = 97;
// bram[21863] = 81;
// bram[21864] = 66;
// bram[21865] = 52;
// bram[21866] = 40;
// bram[21867] = 29;
// bram[21868] = 19;
// bram[21869] = 11;
// bram[21870] = 5;
// bram[21871] = 1;
// bram[21872] = 0;
// bram[21873] = 0;
// bram[21874] = 2;
// bram[21875] = 7;
// bram[21876] = 13;
// bram[21877] = 22;
// bram[21878] = 32;
// bram[21879] = 44;
// bram[21880] = 57;
// bram[21881] = 71;
// bram[21882] = 86;
// bram[21883] = 102;
// bram[21884] = 118;
// bram[21885] = 135;
// bram[21886] = 151;
// bram[21887] = 167;
// bram[21888] = 182;
// bram[21889] = 196;
// bram[21890] = 209;
// bram[21891] = 221;
// bram[21892] = 231;
// bram[21893] = 240;
// bram[21894] = 246;
// bram[21895] = 251;
// bram[21896] = 253;
// bram[21897] = 253;
// bram[21898] = 252;
// bram[21899] = 248;
// bram[21900] = 242;
// bram[21901] = 234;
// bram[21902] = 224;
// bram[21903] = 213;
// bram[21904] = 201;
// bram[21905] = 187;
// bram[21906] = 172;
// bram[21907] = 156;
// bram[21908] = 140;
// bram[21909] = 123;
// bram[21910] = 107;
// bram[21911] = 91;
// bram[21912] = 76;
// bram[21913] = 61;
// bram[21914] = 48;
// bram[21915] = 35;
// bram[21916] = 25;
// bram[21917] = 16;
// bram[21918] = 9;
// bram[21919] = 4;
// bram[21920] = 1;
// bram[21921] = 0;
// bram[21922] = 1;
// bram[21923] = 4;
// bram[21924] = 9;
// bram[21925] = 16;
// bram[21926] = 25;
// bram[21927] = 36;
// bram[21928] = 48;
// bram[21929] = 62;
// bram[21930] = 77;
// bram[21931] = 92;
// bram[21932] = 108;
// bram[21933] = 124;
// bram[21934] = 141;
// bram[21935] = 157;
// bram[21936] = 173;
// bram[21937] = 187;
// bram[21938] = 201;
// bram[21939] = 214;
// bram[21940] = 225;
// bram[21941] = 234;
// bram[21942] = 242;
// bram[21943] = 248;
// bram[21944] = 252;
// bram[21945] = 253;
// bram[21946] = 253;
// bram[21947] = 250;
// bram[21948] = 246;
// bram[21949] = 239;
// bram[21950] = 231;
// bram[21951] = 220;
// bram[21952] = 209;
// bram[21953] = 196;
// bram[21954] = 181;
// bram[21955] = 166;
// bram[21956] = 150;
// bram[21957] = 134;
// bram[21958] = 117;
// bram[21959] = 101;
// bram[21960] = 85;
// bram[21961] = 70;
// bram[21962] = 56;
// bram[21963] = 43;
// bram[21964] = 31;
// bram[21965] = 21;
// bram[21966] = 13;
// bram[21967] = 7;
// bram[21968] = 2;
// bram[21969] = 0;
// bram[21970] = 0;
// bram[21971] = 2;
// bram[21972] = 6;
// bram[21973] = 12;
// bram[21974] = 19;
// bram[21975] = 29;
// bram[21976] = 40;
// bram[21977] = 53;
// bram[21978] = 67;
// bram[21979] = 82;
// bram[21980] = 98;
// bram[21981] = 114;
// bram[21982] = 130;
// bram[21983] = 147;
// bram[21984] = 163;
// bram[21985] = 178;
// bram[21986] = 193;
// bram[21987] = 206;
// bram[21988] = 218;
// bram[21989] = 229;
// bram[21990] = 238;
// bram[21991] = 245;
// bram[21992] = 250;
// bram[21993] = 253;
// bram[21994] = 253;
// bram[21995] = 252;
// bram[21996] = 249;
// bram[21997] = 244;
// bram[21998] = 236;
// bram[21999] = 227;
// bram[22000] = 216;
// bram[22001] = 204;
// bram[22002] = 190;
// bram[22003] = 176;
// bram[22004] = 160;
// bram[22005] = 144;
// bram[22006] = 128;
// bram[22007] = 111;
// bram[22008] = 95;
// bram[22009] = 80;
// bram[22010] = 65;
// bram[22011] = 51;
// bram[22012] = 39;
// bram[22013] = 27;
// bram[22014] = 18;
// bram[22015] = 10;
// bram[22016] = 5;
// bram[22017] = 1;
// bram[22018] = 0;
// bram[22019] = 0;
// bram[22020] = 3;
// bram[22021] = 8;
// bram[22022] = 14;
// bram[22023] = 23;
// bram[22024] = 33;
// bram[22025] = 45;
// bram[22026] = 58;
// bram[22027] = 73;
// bram[22028] = 88;
// bram[22029] = 104;
// bram[22030] = 120;
// bram[22031] = 136;
// bram[22032] = 153;
// bram[22033] = 168;
// bram[22034] = 184;
// bram[22035] = 198;
// bram[22036] = 211;
// bram[22037] = 222;
// bram[22038] = 232;
// bram[22039] = 240;
// bram[22040] = 247;
// bram[22041] = 251;
// bram[22042] = 253;
// bram[22043] = 253;
// bram[22044] = 251;
// bram[22045] = 247;
// bram[22046] = 241;
// bram[22047] = 233;
// bram[22048] = 223;
// bram[22049] = 212;
// bram[22050] = 199;
// bram[22051] = 185;
// bram[22052] = 170;
// bram[22053] = 154;
// bram[22054] = 138;
// bram[22055] = 122;
// bram[22056] = 105;
// bram[22057] = 89;
// bram[22058] = 74;
// bram[22059] = 60;
// bram[22060] = 46;
// bram[22061] = 34;
// bram[22062] = 24;
// bram[22063] = 15;
// bram[22064] = 8;
// bram[22065] = 3;
// bram[22066] = 0;
// bram[22067] = 0;
// bram[22068] = 1;
// bram[22069] = 4;
// bram[22070] = 10;
// bram[22071] = 17;
// bram[22072] = 26;
// bram[22073] = 37;
// bram[22074] = 50;
// bram[22075] = 63;
// bram[22076] = 78;
// bram[22077] = 94;
// bram[22078] = 110;
// bram[22079] = 126;
// bram[22080] = 142;
// bram[22081] = 159;
// bram[22082] = 174;
// bram[22083] = 189;
// bram[22084] = 203;
// bram[22085] = 215;
// bram[22086] = 226;
// bram[22087] = 235;
// bram[22088] = 243;
// bram[22089] = 248;
// bram[22090] = 252;
// bram[22091] = 253;
// bram[22092] = 253;
// bram[22093] = 250;
// bram[22094] = 245;
// bram[22095] = 238;
// bram[22096] = 230;
// bram[22097] = 219;
// bram[22098] = 207;
// bram[22099] = 194;
// bram[22100] = 180;
// bram[22101] = 164;
// bram[22102] = 148;
// bram[22103] = 132;
// bram[22104] = 116;
// bram[22105] = 100;
// bram[22106] = 84;
// bram[22107] = 69;
// bram[22108] = 55;
// bram[22109] = 42;
// bram[22110] = 30;
// bram[22111] = 20;
// bram[22112] = 12;
// bram[22113] = 6;
// bram[22114] = 2;
// bram[22115] = 0;
// bram[22116] = 0;
// bram[22117] = 2;
// bram[22118] = 6;
// bram[22119] = 12;
// bram[22120] = 20;
// bram[22121] = 30;
// bram[22122] = 42;
// bram[22123] = 55;
// bram[22124] = 69;
// bram[22125] = 84;
// bram[22126] = 99;
// bram[22127] = 116;
// bram[22128] = 132;
// bram[22129] = 148;
// bram[22130] = 164;
// bram[22131] = 180;
// bram[22132] = 194;
// bram[22133] = 207;
// bram[22134] = 219;
// bram[22135] = 230;
// bram[22136] = 238;
// bram[22137] = 245;
// bram[22138] = 250;
// bram[22139] = 253;
// bram[22140] = 253;
// bram[22141] = 252;
// bram[22142] = 248;
// bram[22143] = 243;
// bram[22144] = 235;
// bram[22145] = 226;
// bram[22146] = 215;
// bram[22147] = 203;
// bram[22148] = 189;
// bram[22149] = 174;
// bram[22150] = 159;
// bram[22151] = 142;
// bram[22152] = 126;
// bram[22153] = 110;
// bram[22154] = 94;
// bram[22155] = 78;
// bram[22156] = 63;
// bram[22157] = 50;
// bram[22158] = 37;
// bram[22159] = 26;
// bram[22160] = 17;
// bram[22161] = 10;
// bram[22162] = 4;
// bram[22163] = 1;
// bram[22164] = 0;
// bram[22165] = 0;
// bram[22166] = 3;
// bram[22167] = 8;
// bram[22168] = 15;
// bram[22169] = 24;
// bram[22170] = 34;
// bram[22171] = 46;
// bram[22172] = 60;
// bram[22173] = 74;
// bram[22174] = 89;
// bram[22175] = 105;
// bram[22176] = 122;
// bram[22177] = 138;
// bram[22178] = 154;
// bram[22179] = 170;
// bram[22180] = 185;
// bram[22181] = 199;
// bram[22182] = 212;
// bram[22183] = 223;
// bram[22184] = 233;
// bram[22185] = 241;
// bram[22186] = 247;
// bram[22187] = 251;
// bram[22188] = 253;
// bram[22189] = 253;
// bram[22190] = 251;
// bram[22191] = 247;
// bram[22192] = 240;
// bram[22193] = 232;
// bram[22194] = 222;
// bram[22195] = 211;
// bram[22196] = 198;
// bram[22197] = 184;
// bram[22198] = 168;
// bram[22199] = 153;
// bram[22200] = 136;
// bram[22201] = 120;
// bram[22202] = 104;
// bram[22203] = 88;
// bram[22204] = 73;
// bram[22205] = 58;
// bram[22206] = 45;
// bram[22207] = 33;
// bram[22208] = 23;
// bram[22209] = 14;
// bram[22210] = 8;
// bram[22211] = 3;
// bram[22212] = 0;
// bram[22213] = 0;
// bram[22214] = 1;
// bram[22215] = 5;
// bram[22216] = 10;
// bram[22217] = 18;
// bram[22218] = 27;
// bram[22219] = 39;
// bram[22220] = 51;
// bram[22221] = 65;
// bram[22222] = 80;
// bram[22223] = 95;
// bram[22224] = 111;
// bram[22225] = 128;
// bram[22226] = 144;
// bram[22227] = 160;
// bram[22228] = 176;
// bram[22229] = 190;
// bram[22230] = 204;
// bram[22231] = 216;
// bram[22232] = 227;
// bram[22233] = 236;
// bram[22234] = 244;
// bram[22235] = 249;
// bram[22236] = 252;
// bram[22237] = 253;
// bram[22238] = 253;
// bram[22239] = 250;
// bram[22240] = 245;
// bram[22241] = 238;
// bram[22242] = 229;
// bram[22243] = 218;
// bram[22244] = 206;
// bram[22245] = 193;
// bram[22246] = 178;
// bram[22247] = 163;
// bram[22248] = 147;
// bram[22249] = 130;
// bram[22250] = 114;
// bram[22251] = 98;
// bram[22252] = 82;
// bram[22253] = 67;
// bram[22254] = 53;
// bram[22255] = 40;
// bram[22256] = 29;
// bram[22257] = 19;
// bram[22258] = 12;
// bram[22259] = 6;
// bram[22260] = 2;
// bram[22261] = 0;
// bram[22262] = 0;
// bram[22263] = 2;
// bram[22264] = 7;
// bram[22265] = 13;
// bram[22266] = 21;
// bram[22267] = 31;
// bram[22268] = 43;
// bram[22269] = 56;
// bram[22270] = 70;
// bram[22271] = 85;
// bram[22272] = 101;
// bram[22273] = 117;
// bram[22274] = 134;
// bram[22275] = 150;
// bram[22276] = 166;
// bram[22277] = 181;
// bram[22278] = 195;
// bram[22279] = 209;
// bram[22280] = 220;
// bram[22281] = 231;
// bram[22282] = 239;
// bram[22283] = 246;
// bram[22284] = 250;
// bram[22285] = 253;
// bram[22286] = 253;
// bram[22287] = 252;
// bram[22288] = 248;
// bram[22289] = 242;
// bram[22290] = 235;
// bram[22291] = 225;
// bram[22292] = 214;
// bram[22293] = 201;
// bram[22294] = 187;
// bram[22295] = 173;
// bram[22296] = 157;
// bram[22297] = 141;
// bram[22298] = 124;
// bram[22299] = 108;
// bram[22300] = 92;
// bram[22301] = 77;
// bram[22302] = 62;
// bram[22303] = 48;
// bram[22304] = 36;
// bram[22305] = 25;
// bram[22306] = 16;
// bram[22307] = 9;
// bram[22308] = 4;
// bram[22309] = 1;
// bram[22310] = 0;
// bram[22311] = 0;
// bram[22312] = 4;
// bram[22313] = 9;
// bram[22314] = 16;
// bram[22315] = 25;
// bram[22316] = 35;
// bram[22317] = 48;
// bram[22318] = 61;
// bram[22319] = 76;
// bram[22320] = 91;
// bram[22321] = 107;
// bram[22322] = 123;
// bram[22323] = 140;
// bram[22324] = 156;
// bram[22325] = 172;
// bram[22326] = 187;
// bram[22327] = 200;
// bram[22328] = 213;
// bram[22329] = 224;
// bram[22330] = 234;
// bram[22331] = 242;
// bram[22332] = 248;
// bram[22333] = 252;
// bram[22334] = 253;
// bram[22335] = 253;
// bram[22336] = 251;
// bram[22337] = 246;
// bram[22338] = 240;
// bram[22339] = 231;
// bram[22340] = 221;
// bram[22341] = 209;
// bram[22342] = 196;
// bram[22343] = 182;
// bram[22344] = 167;
// bram[22345] = 151;
// bram[22346] = 135;
// bram[22347] = 118;
// bram[22348] = 102;
// bram[22349] = 86;
// bram[22350] = 71;
// bram[22351] = 57;
// bram[22352] = 44;
// bram[22353] = 32;
// bram[22354] = 22;
// bram[22355] = 13;
// bram[22356] = 7;
// bram[22357] = 2;
// bram[22358] = 0;
// bram[22359] = 0;
// bram[22360] = 1;
// bram[22361] = 5;
// bram[22362] = 11;
// bram[22363] = 19;
// bram[22364] = 29;
// bram[22365] = 40;
// bram[22366] = 52;
// bram[22367] = 66;
// bram[22368] = 81;
// bram[22369] = 97;
// bram[22370] = 113;
// bram[22371] = 129;
// bram[22372] = 146;
// bram[22373] = 162;
// bram[22374] = 177;
// bram[22375] = 192;
// bram[22376] = 205;
// bram[22377] = 217;
// bram[22378] = 228;
// bram[22379] = 237;
// bram[22380] = 244;
// bram[22381] = 249;
// bram[22382] = 252;
// bram[22383] = 253;
// bram[22384] = 252;
// bram[22385] = 249;
// bram[22386] = 244;
// bram[22387] = 237;
// bram[22388] = 228;
// bram[22389] = 217;
// bram[22390] = 205;
// bram[22391] = 191;
// bram[22392] = 177;
// bram[22393] = 161;
// bram[22394] = 145;
// bram[22395] = 129;
// bram[22396] = 112;
// bram[22397] = 96;
// bram[22398] = 81;
// bram[22399] = 66;
// bram[22400] = 52;
// bram[22401] = 39;
// bram[22402] = 28;
// bram[22403] = 19;
// bram[22404] = 11;
// bram[22405] = 5;
// bram[22406] = 1;
// bram[22407] = 0;
// bram[22408] = 0;
// bram[22409] = 3;
// bram[22410] = 7;
// bram[22411] = 14;
// bram[22412] = 22;
// bram[22413] = 32;
// bram[22414] = 44;
// bram[22415] = 57;
// bram[22416] = 72;
// bram[22417] = 87;
// bram[22418] = 103;
// bram[22419] = 119;
// bram[22420] = 135;
// bram[22421] = 152;
// bram[22422] = 168;
// bram[22423] = 183;
// bram[22424] = 197;
// bram[22425] = 210;
// bram[22426] = 222;
// bram[22427] = 232;
// bram[22428] = 240;
// bram[22429] = 246;
// bram[22430] = 251;
// bram[22431] = 253;
// bram[22432] = 253;
// bram[22433] = 251;
// bram[22434] = 247;
// bram[22435] = 242;
// bram[22436] = 234;
// bram[22437] = 224;
// bram[22438] = 213;
// bram[22439] = 200;
// bram[22440] = 186;
// bram[22441] = 171;
// bram[22442] = 155;
// bram[22443] = 139;
// bram[22444] = 123;
// bram[22445] = 106;
// bram[22446] = 90;
// bram[22447] = 75;
// bram[22448] = 60;
// bram[22449] = 47;
// bram[22450] = 35;
// bram[22451] = 24;
// bram[22452] = 15;
// bram[22453] = 8;
// bram[22454] = 3;
// bram[22455] = 0;
// bram[22456] = 0;
// bram[22457] = 1;
// bram[22458] = 4;
// bram[22459] = 9;
// bram[22460] = 17;
// bram[22461] = 26;
// bram[22462] = 37;
// bram[22463] = 49;
// bram[22464] = 63;
// bram[22465] = 77;
// bram[22466] = 93;
// bram[22467] = 109;
// bram[22468] = 125;
// bram[22469] = 141;
// bram[22470] = 158;
// bram[22471] = 173;
// bram[22472] = 188;
// bram[22473] = 202;
// bram[22474] = 214;
// bram[22475] = 225;
// bram[22476] = 235;
// bram[22477] = 243;
// bram[22478] = 248;
// bram[22479] = 252;
// bram[22480] = 253;
// bram[22481] = 253;
// bram[22482] = 250;
// bram[22483] = 246;
// bram[22484] = 239;
// bram[22485] = 230;
// bram[22486] = 220;
// bram[22487] = 208;
// bram[22488] = 195;
// bram[22489] = 181;
// bram[22490] = 165;
// bram[22491] = 149;
// bram[22492] = 133;
// bram[22493] = 117;
// bram[22494] = 100;
// bram[22495] = 85;
// bram[22496] = 70;
// bram[22497] = 55;
// bram[22498] = 42;
// bram[22499] = 31;
// bram[22500] = 21;
// bram[22501] = 13;
// bram[22502] = 6;
// bram[22503] = 2;
// bram[22504] = 0;
// bram[22505] = 0;
// bram[22506] = 2;
// bram[22507] = 6;
// bram[22508] = 12;
// bram[22509] = 20;
// bram[22510] = 30;
// bram[22511] = 41;
// bram[22512] = 54;
// bram[22513] = 68;
// bram[22514] = 83;
// bram[22515] = 99;
// bram[22516] = 115;
// bram[22517] = 131;
// bram[22518] = 147;
// bram[22519] = 163;
// bram[22520] = 179;
// bram[22521] = 193;
// bram[22522] = 207;
// bram[22523] = 219;
// bram[22524] = 229;
// bram[22525] = 238;
// bram[22526] = 245;
// bram[22527] = 250;
// bram[22528] = 253;
// bram[22529] = 253;
// bram[22530] = 252;
// bram[22531] = 249;
// bram[22532] = 243;
// bram[22533] = 236;
// bram[22534] = 227;
// bram[22535] = 216;
// bram[22536] = 203;
// bram[22537] = 190;
// bram[22538] = 175;
// bram[22539] = 159;
// bram[22540] = 143;
// bram[22541] = 127;
// bram[22542] = 111;
// bram[22543] = 95;
// bram[22544] = 79;
// bram[22545] = 64;
// bram[22546] = 50;
// bram[22547] = 38;
// bram[22548] = 27;
// bram[22549] = 18;
// bram[22550] = 10;
// bram[22551] = 5;
// bram[22552] = 1;
// bram[22553] = 0;
// bram[22554] = 0;
// bram[22555] = 3;
// bram[22556] = 8;
// bram[22557] = 15;
// bram[22558] = 23;
// bram[22559] = 34;
// bram[22560] = 46;
// bram[22561] = 59;
// bram[22562] = 73;
// bram[22563] = 89;
// bram[22564] = 104;
// bram[22565] = 121;
// bram[22566] = 137;
// bram[22567] = 153;
// bram[22568] = 169;
// bram[22569] = 184;
// bram[22570] = 198;
// bram[22571] = 211;
// bram[22572] = 223;
// bram[22573] = 233;
// bram[22574] = 241;
// bram[22575] = 247;
// bram[22576] = 251;
// bram[22577] = 253;
// bram[22578] = 253;
// bram[22579] = 251;
// bram[22580] = 247;
// bram[22581] = 241;
// bram[22582] = 233;
// bram[22583] = 223;
// bram[22584] = 211;
// bram[22585] = 199;
// bram[22586] = 184;
// bram[22587] = 169;
// bram[22588] = 154;
// bram[22589] = 137;
// bram[22590] = 121;
// bram[22591] = 105;
// bram[22592] = 89;
// bram[22593] = 73;
// bram[22594] = 59;
// bram[22595] = 46;
// bram[22596] = 34;
// bram[22597] = 23;
// bram[22598] = 15;
// bram[22599] = 8;
// bram[22600] = 3;
// bram[22601] = 0;
// bram[22602] = 0;
// bram[22603] = 1;
// bram[22604] = 4;
// bram[22605] = 10;
// bram[22606] = 18;
// bram[22607] = 27;
// bram[22608] = 38;
// bram[22609] = 50;
// bram[22610] = 64;
// bram[22611] = 79;
// bram[22612] = 94;
// bram[22613] = 110;
// bram[22614] = 127;
// bram[22615] = 143;
// bram[22616] = 159;
// bram[22617] = 175;
// bram[22618] = 190;
// bram[22619] = 203;
// bram[22620] = 216;
// bram[22621] = 227;
// bram[22622] = 236;
// bram[22623] = 243;
// bram[22624] = 249;
// bram[22625] = 252;
// bram[22626] = 253;
// bram[22627] = 253;
// bram[22628] = 250;
// bram[22629] = 245;
// bram[22630] = 238;
// bram[22631] = 229;
// bram[22632] = 219;
// bram[22633] = 207;
// bram[22634] = 193;
// bram[22635] = 179;
// bram[22636] = 164;
// bram[22637] = 148;
// bram[22638] = 131;
// bram[22639] = 115;
// bram[22640] = 99;
// bram[22641] = 83;
// bram[22642] = 68;
// bram[22643] = 54;
// bram[22644] = 41;
// bram[22645] = 30;
// bram[22646] = 20;
// bram[22647] = 12;
// bram[22648] = 6;
// bram[22649] = 2;
// bram[22650] = 0;
// bram[22651] = 0;
// bram[22652] = 2;
// bram[22653] = 6;
// bram[22654] = 13;
// bram[22655] = 21;
// bram[22656] = 31;
// bram[22657] = 42;
// bram[22658] = 55;
// bram[22659] = 69;
// bram[22660] = 84;
// bram[22661] = 100;
// bram[22662] = 116;
// bram[22663] = 133;
// bram[22664] = 149;
// bram[22665] = 165;
// bram[22666] = 180;
// bram[22667] = 195;
// bram[22668] = 208;
// bram[22669] = 220;
// bram[22670] = 230;
// bram[22671] = 239;
// bram[22672] = 245;
// bram[22673] = 250;
// bram[22674] = 253;
// bram[22675] = 253;
// bram[22676] = 252;
// bram[22677] = 248;
// bram[22678] = 243;
// bram[22679] = 235;
// bram[22680] = 226;
// bram[22681] = 215;
// bram[22682] = 202;
// bram[22683] = 188;
// bram[22684] = 173;
// bram[22685] = 158;
// bram[22686] = 142;
// bram[22687] = 125;
// bram[22688] = 109;
// bram[22689] = 93;
// bram[22690] = 77;
// bram[22691] = 63;
// bram[22692] = 49;
// bram[22693] = 37;
// bram[22694] = 26;
// bram[22695] = 17;
// bram[22696] = 9;
// bram[22697] = 4;
// bram[22698] = 1;
// bram[22699] = 0;
// bram[22700] = 0;
// bram[22701] = 3;
// bram[22702] = 8;
// bram[22703] = 15;
// bram[22704] = 24;
// bram[22705] = 35;
// bram[22706] = 47;
// bram[22707] = 60;
// bram[22708] = 75;
// bram[22709] = 90;
// bram[22710] = 106;
// bram[22711] = 122;
// bram[22712] = 139;
// bram[22713] = 155;
// bram[22714] = 171;
// bram[22715] = 186;
// bram[22716] = 200;
// bram[22717] = 212;
// bram[22718] = 224;
// bram[22719] = 233;
// bram[22720] = 241;
// bram[22721] = 247;
// bram[22722] = 251;
// bram[22723] = 253;
// bram[22724] = 253;
// bram[22725] = 251;
// bram[22726] = 246;
// bram[22727] = 240;
// bram[22728] = 232;
// bram[22729] = 222;
// bram[22730] = 210;
// bram[22731] = 197;
// bram[22732] = 183;
// bram[22733] = 168;
// bram[22734] = 152;
// bram[22735] = 136;
// bram[22736] = 119;
// bram[22737] = 103;
// bram[22738] = 87;
// bram[22739] = 72;
// bram[22740] = 58;
// bram[22741] = 44;
// bram[22742] = 33;
// bram[22743] = 22;
// bram[22744] = 14;
// bram[22745] = 7;
// bram[22746] = 3;
// bram[22747] = 0;
// bram[22748] = 0;
// bram[22749] = 1;
// bram[22750] = 5;
// bram[22751] = 11;
// bram[22752] = 18;
// bram[22753] = 28;
// bram[22754] = 39;
// bram[22755] = 52;
// bram[22756] = 65;
// bram[22757] = 80;
// bram[22758] = 96;
// bram[22759] = 112;
// bram[22760] = 128;
// bram[22761] = 145;
// bram[22762] = 161;
// bram[22763] = 176;
// bram[22764] = 191;
// bram[22765] = 205;
// bram[22766] = 217;
// bram[22767] = 228;
// bram[22768] = 237;
// bram[22769] = 244;
// bram[22770] = 249;
// bram[22771] = 252;
// bram[22772] = 253;
// bram[22773] = 253;
// bram[22774] = 249;
// bram[22775] = 244;
// bram[22776] = 237;
// bram[22777] = 228;
// bram[22778] = 218;
// bram[22779] = 205;
// bram[22780] = 192;
// bram[22781] = 177;
// bram[22782] = 162;
// bram[22783] = 146;
// bram[22784] = 130;
// bram[22785] = 113;
// bram[22786] = 97;
// bram[22787] = 81;
// bram[22788] = 67;
// bram[22789] = 53;
// bram[22790] = 40;
// bram[22791] = 29;
// bram[22792] = 19;
// bram[22793] = 11;
// bram[22794] = 5;
// bram[22795] = 1;
// bram[22796] = 0;
// bram[22797] = 0;
// bram[22798] = 2;
// bram[22799] = 7;
// bram[22800] = 13;
// bram[22801] = 22;
// bram[22802] = 32;
// bram[22803] = 44;
// bram[22804] = 57;
// bram[22805] = 71;
// bram[22806] = 86;
// bram[22807] = 102;
// bram[22808] = 118;
// bram[22809] = 135;
// bram[22810] = 151;
// bram[22811] = 167;
// bram[22812] = 182;
// bram[22813] = 196;
// bram[22814] = 209;
// bram[22815] = 221;
// bram[22816] = 231;
// bram[22817] = 239;
// bram[22818] = 246;
// bram[22819] = 251;
// bram[22820] = 253;
// bram[22821] = 253;
// bram[22822] = 252;
// bram[22823] = 248;
// bram[22824] = 242;
// bram[22825] = 234;
// bram[22826] = 225;
// bram[22827] = 213;
// bram[22828] = 201;
// bram[22829] = 187;
// bram[22830] = 172;
// bram[22831] = 156;
// bram[22832] = 140;
// bram[22833] = 124;
// bram[22834] = 107;
// bram[22835] = 91;
// bram[22836] = 76;
// bram[22837] = 61;
// bram[22838] = 48;
// bram[22839] = 36;
// bram[22840] = 25;
// bram[22841] = 16;
// bram[22842] = 9;
// bram[22843] = 4;
// bram[22844] = 1;
// bram[22845] = 0;
// bram[22846] = 1;
// bram[22847] = 4;
// bram[22848] = 9;
// bram[22849] = 16;
// bram[22850] = 25;
// bram[22851] = 36;
// bram[22852] = 48;
// bram[22853] = 62;
// bram[22854] = 76;
// bram[22855] = 92;
// bram[22856] = 108;
// bram[22857] = 124;
// bram[22858] = 141;
// bram[22859] = 157;
// bram[22860] = 172;
// bram[22861] = 187;
// bram[22862] = 201;
// bram[22863] = 214;
// bram[22864] = 225;
// bram[22865] = 234;
// bram[22866] = 242;
// bram[22867] = 248;
// bram[22868] = 252;
// bram[22869] = 253;
// bram[22870] = 253;
// bram[22871] = 250;
// bram[22872] = 246;
// bram[22873] = 239;
// bram[22874] = 231;
// bram[22875] = 221;
// bram[22876] = 209;
// bram[22877] = 196;
// bram[22878] = 181;
// bram[22879] = 166;
// bram[22880] = 150;
// bram[22881] = 134;
// bram[22882] = 118;
// bram[22883] = 101;
// bram[22884] = 86;
// bram[22885] = 70;
// bram[22886] = 56;
// bram[22887] = 43;
// bram[22888] = 32;
// bram[22889] = 21;
// bram[22890] = 13;
// bram[22891] = 7;
// bram[22892] = 2;
// bram[22893] = 0;
// bram[22894] = 0;
// bram[22895] = 2;
// bram[22896] = 5;
// bram[22897] = 11;
// bram[22898] = 19;
// bram[22899] = 29;
// bram[22900] = 40;
// bram[22901] = 53;
// bram[22902] = 67;
// bram[22903] = 82;
// bram[22904] = 98;
// bram[22905] = 114;
// bram[22906] = 130;
// bram[22907] = 147;
// bram[22908] = 163;
// bram[22909] = 178;
// bram[22910] = 192;
// bram[22911] = 206;
// bram[22912] = 218;
// bram[22913] = 229;
// bram[22914] = 237;
// bram[22915] = 244;
// bram[22916] = 250;
// bram[22917] = 253;
// bram[22918] = 253;
// bram[22919] = 252;
// bram[22920] = 249;
// bram[22921] = 244;
// bram[22922] = 236;
// bram[22923] = 227;
// bram[22924] = 216;
// bram[22925] = 204;
// bram[22926] = 191;
// bram[22927] = 176;
// bram[22928] = 160;
// bram[22929] = 144;
// bram[22930] = 128;
// bram[22931] = 112;
// bram[22932] = 95;
// bram[22933] = 80;
// bram[22934] = 65;
// bram[22935] = 51;
// bram[22936] = 39;
// bram[22937] = 28;
// bram[22938] = 18;
// bram[22939] = 11;
// bram[22940] = 5;
// bram[22941] = 1;
// bram[22942] = 0;
// bram[22943] = 0;
// bram[22944] = 3;
// bram[22945] = 7;
// bram[22946] = 14;
// bram[22947] = 23;
// bram[22948] = 33;
// bram[22949] = 45;
// bram[22950] = 58;
// bram[22951] = 72;
// bram[22952] = 88;
// bram[22953] = 104;
// bram[22954] = 120;
// bram[22955] = 136;
// bram[22956] = 152;
// bram[22957] = 168;
// bram[22958] = 183;
// bram[22959] = 198;
// bram[22960] = 210;
// bram[22961] = 222;
// bram[22962] = 232;
// bram[22963] = 240;
// bram[22964] = 247;
// bram[22965] = 251;
// bram[22966] = 253;
// bram[22967] = 253;
// bram[22968] = 251;
// bram[22969] = 247;
// bram[22970] = 241;
// bram[22971] = 233;
// bram[22972] = 223;
// bram[22973] = 212;
// bram[22974] = 199;
// bram[22975] = 185;
// bram[22976] = 170;
// bram[22977] = 155;
// bram[22978] = 138;
// bram[22979] = 122;
// bram[22980] = 106;
// bram[22981] = 90;
// bram[22982] = 74;
// bram[22983] = 60;
// bram[22984] = 46;
// bram[22985] = 34;
// bram[22986] = 24;
// bram[22987] = 15;
// bram[22988] = 8;
// bram[22989] = 3;
// bram[22990] = 0;
// bram[22991] = 0;
// bram[22992] = 1;
// bram[22993] = 4;
// bram[22994] = 10;
// bram[22995] = 17;
// bram[22996] = 26;
// bram[22997] = 37;
// bram[22998] = 50;
// bram[22999] = 63;
// bram[23000] = 78;
// bram[23001] = 93;
// bram[23002] = 109;
// bram[23003] = 126;
// bram[23004] = 142;
// bram[23005] = 158;
// bram[23006] = 174;
// bram[23007] = 189;
// bram[23008] = 202;
// bram[23009] = 215;
// bram[23010] = 226;
// bram[23011] = 235;
// bram[23012] = 243;
// bram[23013] = 248;
// bram[23014] = 252;
// bram[23015] = 253;
// bram[23016] = 253;
// bram[23017] = 250;
// bram[23018] = 245;
// bram[23019] = 238;
// bram[23020] = 230;
// bram[23021] = 219;
// bram[23022] = 208;
// bram[23023] = 194;
// bram[23024] = 180;
// bram[23025] = 165;
// bram[23026] = 149;
// bram[23027] = 132;
// bram[23028] = 116;
// bram[23029] = 100;
// bram[23030] = 84;
// bram[23031] = 69;
// bram[23032] = 55;
// bram[23033] = 42;
// bram[23034] = 30;
// bram[23035] = 20;
// bram[23036] = 12;
// bram[23037] = 6;
// bram[23038] = 2;
// bram[23039] = 0;
// bram[23040] = 0;
// bram[23041] = 2;
// bram[23042] = 6;
// bram[23043] = 12;
// bram[23044] = 20;
// bram[23045] = 30;
// bram[23046] = 42;
// bram[23047] = 54;
// bram[23048] = 68;
// bram[23049] = 84;
// bram[23050] = 99;
// bram[23051] = 115;
// bram[23052] = 132;
// bram[23053] = 148;
// bram[23054] = 164;
// bram[23055] = 179;
// bram[23056] = 194;
// bram[23057] = 207;
// bram[23058] = 219;
// bram[23059] = 230;
// bram[23060] = 238;
// bram[23061] = 245;
// bram[23062] = 250;
// bram[23063] = 253;
// bram[23064] = 253;
// bram[23065] = 252;
// bram[23066] = 249;
// bram[23067] = 243;
// bram[23068] = 236;
// bram[23069] = 226;
// bram[23070] = 215;
// bram[23071] = 203;
// bram[23072] = 189;
// bram[23073] = 174;
// bram[23074] = 159;
// bram[23075] = 143;
// bram[23076] = 126;
// bram[23077] = 110;
// bram[23078] = 94;
// bram[23079] = 78;
// bram[23080] = 64;
// bram[23081] = 50;
// bram[23082] = 37;
// bram[23083] = 27;
// bram[23084] = 17;
// bram[23085] = 10;
// bram[23086] = 4;
// bram[23087] = 1;
// bram[23088] = 0;
// bram[23089] = 0;
// bram[23090] = 3;
// bram[23091] = 8;
// bram[23092] = 15;
// bram[23093] = 24;
// bram[23094] = 34;
// bram[23095] = 46;
// bram[23096] = 59;
// bram[23097] = 74;
// bram[23098] = 89;
// bram[23099] = 105;
// bram[23100] = 122;
// bram[23101] = 138;
// bram[23102] = 154;
// bram[23103] = 170;
// bram[23104] = 185;
// bram[23105] = 199;
// bram[23106] = 212;
// bram[23107] = 223;
// bram[23108] = 233;
// bram[23109] = 241;
// bram[23110] = 247;
// bram[23111] = 251;
// bram[23112] = 253;
// bram[23113] = 253;
// bram[23114] = 251;
// bram[23115] = 247;
// bram[23116] = 240;
// bram[23117] = 232;
// bram[23118] = 222;
// bram[23119] = 211;
// bram[23120] = 198;
// bram[23121] = 184;
// bram[23122] = 169;
// bram[23123] = 153;
// bram[23124] = 137;
// bram[23125] = 120;
// bram[23126] = 104;
// bram[23127] = 88;
// bram[23128] = 73;
// bram[23129] = 58;
// bram[23130] = 45;
// bram[23131] = 33;
// bram[23132] = 23;
// bram[23133] = 14;
// bram[23134] = 8;
// bram[23135] = 3;
// bram[23136] = 0;
// bram[23137] = 0;
// bram[23138] = 1;
// bram[23139] = 5;
// bram[23140] = 10;
// bram[23141] = 18;
// bram[23142] = 27;
// bram[23143] = 38;
// bram[23144] = 51;
// bram[23145] = 65;
// bram[23146] = 79;
// bram[23147] = 95;
// bram[23148] = 111;
// bram[23149] = 128;
// bram[23150] = 144;
// bram[23151] = 160;
// bram[23152] = 175;
// bram[23153] = 190;
// bram[23154] = 204;
// bram[23155] = 216;
// bram[23156] = 227;
// bram[23157] = 236;
// bram[23158] = 243;
// bram[23159] = 249;
// bram[23160] = 252;
// bram[23161] = 253;
// bram[23162] = 253;
// bram[23163] = 250;
// bram[23164] = 245;
// bram[23165] = 238;
// bram[23166] = 229;
// bram[23167] = 218;
// bram[23168] = 206;
// bram[23169] = 193;
// bram[23170] = 178;
// bram[23171] = 163;
// bram[23172] = 147;
// bram[23173] = 131;
// bram[23174] = 114;
// bram[23175] = 98;
// bram[23176] = 82;
// bram[23177] = 67;
// bram[23178] = 53;
// bram[23179] = 41;
// bram[23180] = 29;
// bram[23181] = 20;
// bram[23182] = 12;
// bram[23183] = 6;
// bram[23184] = 2;
// bram[23185] = 0;
// bram[23186] = 0;
// bram[23187] = 2;
// bram[23188] = 7;
// bram[23189] = 13;
// bram[23190] = 21;
// bram[23191] = 31;
// bram[23192] = 43;
// bram[23193] = 56;
// bram[23194] = 70;
// bram[23195] = 85;
// bram[23196] = 101;
// bram[23197] = 117;
// bram[23198] = 134;
// bram[23199] = 150;
// bram[23200] = 166;
// bram[23201] = 181;
// bram[23202] = 195;
// bram[23203] = 208;
// bram[23204] = 220;
// bram[23205] = 231;
// bram[23206] = 239;
// bram[23207] = 246;
// bram[23208] = 250;
// bram[23209] = 253;
// bram[23210] = 253;
// bram[23211] = 252;
// bram[23212] = 248;
// bram[23213] = 242;
// bram[23214] = 235;
// bram[23215] = 225;
// bram[23216] = 214;
// bram[23217] = 201;
// bram[23218] = 188;
// bram[23219] = 173;
// bram[23220] = 157;
// bram[23221] = 141;
// bram[23222] = 125;
// bram[23223] = 108;
// bram[23224] = 92;
// bram[23225] = 77;
// bram[23226] = 62;
// bram[23227] = 49;
// bram[23228] = 36;
// bram[23229] = 26;
// bram[23230] = 16;
// bram[23231] = 9;
// bram[23232] = 4;
// bram[23233] = 1;
// bram[23234] = 0;
// bram[23235] = 0;
// bram[23236] = 4;
// bram[23237] = 9;
// bram[23238] = 16;
// bram[23239] = 25;
// bram[23240] = 35;
// bram[23241] = 47;
// bram[23242] = 61;
// bram[23243] = 75;
// bram[23244] = 91;
// bram[23245] = 107;
// bram[23246] = 123;
// bram[23247] = 140;
// bram[23248] = 156;
// bram[23249] = 171;
// bram[23250] = 186;
// bram[23251] = 200;
// bram[23252] = 213;
// bram[23253] = 224;
// bram[23254] = 234;
// bram[23255] = 242;
// bram[23256] = 248;
// bram[23257] = 252;
// bram[23258] = 253;
// bram[23259] = 253;
// bram[23260] = 251;
// bram[23261] = 246;
// bram[23262] = 240;
// bram[23263] = 231;
// bram[23264] = 221;
// bram[23265] = 210;
// bram[23266] = 196;
// bram[23267] = 182;
// bram[23268] = 167;
// bram[23269] = 151;
// bram[23270] = 135;
// bram[23271] = 119;
// bram[23272] = 102;
// bram[23273] = 86;
// bram[23274] = 71;
// bram[23275] = 57;
// bram[23276] = 44;
// bram[23277] = 32;
// bram[23278] = 22;
// bram[23279] = 14;
// bram[23280] = 7;
// bram[23281] = 2;
// bram[23282] = 0;
// bram[23283] = 0;
// bram[23284] = 1;
// bram[23285] = 5;
// bram[23286] = 11;
// bram[23287] = 19;
// bram[23288] = 28;
// bram[23289] = 40;
// bram[23290] = 52;
// bram[23291] = 66;
// bram[23292] = 81;
// bram[23293] = 97;
// bram[23294] = 113;
// bram[23295] = 129;
// bram[23296] = 146;
// bram[23297] = 162;
// bram[23298] = 177;
// bram[23299] = 192;
// bram[23300] = 205;
// bram[23301] = 217;
// bram[23302] = 228;
// bram[23303] = 237;
// bram[23304] = 244;
// bram[23305] = 249;
// bram[23306] = 252;
// bram[23307] = 253;
// bram[23308] = 252;
// bram[23309] = 249;
// bram[23310] = 244;
// bram[23311] = 237;
// bram[23312] = 228;
// bram[23313] = 217;
// bram[23314] = 205;
// bram[23315] = 191;
// bram[23316] = 177;
// bram[23317] = 161;
// bram[23318] = 145;
// bram[23319] = 129;
// bram[23320] = 113;
// bram[23321] = 96;
// bram[23322] = 81;
// bram[23323] = 66;
// bram[23324] = 52;
// bram[23325] = 39;
// bram[23326] = 28;
// bram[23327] = 19;
// bram[23328] = 11;
// bram[23329] = 5;
// bram[23330] = 1;
// bram[23331] = 0;
// bram[23332] = 0;
// bram[23333] = 3;
// bram[23334] = 7;
// bram[23335] = 14;
// bram[23336] = 22;
// bram[23337] = 32;
// bram[23338] = 44;
// bram[23339] = 57;
// bram[23340] = 72;
// bram[23341] = 87;
// bram[23342] = 103;
// bram[23343] = 119;
// bram[23344] = 135;
// bram[23345] = 152;
// bram[23346] = 167;
// bram[23347] = 183;
// bram[23348] = 197;
// bram[23349] = 210;
// bram[23350] = 221;
// bram[23351] = 232;
// bram[23352] = 240;
// bram[23353] = 246;
// bram[23354] = 251;
// bram[23355] = 253;
// bram[23356] = 253;
// bram[23357] = 251;
// bram[23358] = 248;
// bram[23359] = 242;
// bram[23360] = 234;
// bram[23361] = 224;
// bram[23362] = 213;
// bram[23363] = 200;
// bram[23364] = 186;
// bram[23365] = 171;
// bram[23366] = 155;
// bram[23367] = 139;
// bram[23368] = 123;
// bram[23369] = 107;
// bram[23370] = 91;
// bram[23371] = 75;
// bram[23372] = 61;
// bram[23373] = 47;
// bram[23374] = 35;
// bram[23375] = 24;
// bram[23376] = 16;
// bram[23377] = 9;
// bram[23378] = 3;
// bram[23379] = 0;
// bram[23380] = 0;
// bram[23381] = 1;
// bram[23382] = 4;
// bram[23383] = 9;
// bram[23384] = 17;
// bram[23385] = 26;
// bram[23386] = 36;
// bram[23387] = 49;
// bram[23388] = 62;
// bram[23389] = 77;
// bram[23390] = 93;
// bram[23391] = 109;
// bram[23392] = 125;
// bram[23393] = 141;
// bram[23394] = 157;
// bram[23395] = 173;
// bram[23396] = 188;
// bram[23397] = 202;
// bram[23398] = 214;
// bram[23399] = 225;
// bram[23400] = 235;
// bram[23401] = 242;
// bram[23402] = 248;
// bram[23403] = 252;
// bram[23404] = 253;
// bram[23405] = 253;
// bram[23406] = 250;
// bram[23407] = 246;
// bram[23408] = 239;
// bram[23409] = 230;
// bram[23410] = 220;
// bram[23411] = 208;
// bram[23412] = 195;
// bram[23413] = 181;
// bram[23414] = 165;
// bram[23415] = 150;
// bram[23416] = 133;
// bram[23417] = 117;
// bram[23418] = 101;
// bram[23419] = 85;
// bram[23420] = 70;
// bram[23421] = 56;
// bram[23422] = 43;
// bram[23423] = 31;
// bram[23424] = 21;
// bram[23425] = 13;
// bram[23426] = 6;
// bram[23427] = 2;
// bram[23428] = 0;
// bram[23429] = 0;
// bram[23430] = 2;
// bram[23431] = 6;
// bram[23432] = 12;
// bram[23433] = 20;
// bram[23434] = 29;
// bram[23435] = 41;
// bram[23436] = 54;
// bram[23437] = 68;
// bram[23438] = 83;
// bram[23439] = 98;
// bram[23440] = 115;
// bram[23441] = 131;
// bram[23442] = 147;
// bram[23443] = 163;
// bram[23444] = 179;
// bram[23445] = 193;
// bram[23446] = 206;
// bram[23447] = 218;
// bram[23448] = 229;
// bram[23449] = 238;
// bram[23450] = 245;
// bram[23451] = 250;
// bram[23452] = 253;
// bram[23453] = 253;
// bram[23454] = 252;
// bram[23455] = 249;
// bram[23456] = 243;
// bram[23457] = 236;
// bram[23458] = 227;
// bram[23459] = 216;
// bram[23460] = 204;
// bram[23461] = 190;
// bram[23462] = 175;
// bram[23463] = 160;
// bram[23464] = 144;
// bram[23465] = 127;
// bram[23466] = 111;
// bram[23467] = 95;
// bram[23468] = 79;
// bram[23469] = 64;
// bram[23470] = 51;
// bram[23471] = 38;
// bram[23472] = 27;
// bram[23473] = 18;
// bram[23474] = 10;
// bram[23475] = 5;
// bram[23476] = 1;
// bram[23477] = 0;
// bram[23478] = 0;
// bram[23479] = 3;
// bram[23480] = 8;
// bram[23481] = 14;
// bram[23482] = 23;
// bram[23483] = 33;
// bram[23484] = 45;
// bram[23485] = 59;
// bram[23486] = 73;
// bram[23487] = 88;
// bram[23488] = 104;
// bram[23489] = 121;
// bram[23490] = 137;
// bram[23491] = 153;
// bram[23492] = 169;
// bram[23493] = 184;
// bram[23494] = 198;
// bram[23495] = 211;
// bram[23496] = 223;
// bram[23497] = 232;
// bram[23498] = 241;
// bram[23499] = 247;
// bram[23500] = 251;
// bram[23501] = 253;
// bram[23502] = 253;
// bram[23503] = 251;
// bram[23504] = 247;
// bram[23505] = 241;
// bram[23506] = 233;
// bram[23507] = 223;
// bram[23508] = 212;
// bram[23509] = 199;
// bram[23510] = 185;
// bram[23511] = 170;
// bram[23512] = 154;
// bram[23513] = 138;
// bram[23514] = 121;
// bram[23515] = 105;
// bram[23516] = 89;
// bram[23517] = 74;
// bram[23518] = 59;
// bram[23519] = 46;
// bram[23520] = 34;
// bram[23521] = 23;
// bram[23522] = 15;
// bram[23523] = 8;
// bram[23524] = 3;
// bram[23525] = 0;
// bram[23526] = 0;
// bram[23527] = 1;
// bram[23528] = 4;
// bram[23529] = 10;
// bram[23530] = 17;
// bram[23531] = 27;
// bram[23532] = 38;
// bram[23533] = 50;
// bram[23534] = 64;
// bram[23535] = 79;
// bram[23536] = 94;
// bram[23537] = 110;
// bram[23538] = 127;
// bram[23539] = 143;
// bram[23540] = 159;
// bram[23541] = 175;
// bram[23542] = 189;
// bram[23543] = 203;
// bram[23544] = 215;
// bram[23545] = 226;
// bram[23546] = 236;
// bram[23547] = 243;
// bram[23548] = 249;
// bram[23549] = 252;
// bram[23550] = 253;
// bram[23551] = 253;
// bram[23552] = 250;
// bram[23553] = 245;
// bram[23554] = 238;
// bram[23555] = 229;
// bram[23556] = 219;
// bram[23557] = 207;
// bram[23558] = 194;
// bram[23559] = 179;
// bram[23560] = 164;
// bram[23561] = 148;
// bram[23562] = 132;
// bram[23563] = 115;
// bram[23564] = 99;
// bram[23565] = 83;
// bram[23566] = 68;
// bram[23567] = 54;
// bram[23568] = 41;
// bram[23569] = 30;
// bram[23570] = 20;
// bram[23571] = 12;
// bram[23572] = 6;
// bram[23573] = 2;
// bram[23574] = 0;
// bram[23575] = 0;
// bram[23576] = 2;
// bram[23577] = 6;
// bram[23578] = 12;
// bram[23579] = 21;
// bram[23580] = 31;
// bram[23581] = 42;
// bram[23582] = 55;
// bram[23583] = 69;
// bram[23584] = 84;
// bram[23585] = 100;
// bram[23586] = 116;
// bram[23587] = 133;
// bram[23588] = 149;
// bram[23589] = 165;
// bram[23590] = 180;
// bram[23591] = 195;
// bram[23592] = 208;
// bram[23593] = 220;
// bram[23594] = 230;
// bram[23595] = 239;
// bram[23596] = 245;
// bram[23597] = 250;
// bram[23598] = 253;
// bram[23599] = 253;
// bram[23600] = 252;
// bram[23601] = 248;
// bram[23602] = 243;
// bram[23603] = 235;
// bram[23604] = 226;
// bram[23605] = 215;
// bram[23606] = 202;
// bram[23607] = 188;
// bram[23608] = 174;
// bram[23609] = 158;
// bram[23610] = 142;
// bram[23611] = 126;
// bram[23612] = 109;
// bram[23613] = 93;
// bram[23614] = 78;
// bram[23615] = 63;
// bram[23616] = 49;
// bram[23617] = 37;
// bram[23618] = 26;
// bram[23619] = 17;
// bram[23620] = 10;
// bram[23621] = 4;
// bram[23622] = 1;
// bram[23623] = 0;
// bram[23624] = 0;
// bram[23625] = 3;
// bram[23626] = 8;
// bram[23627] = 15;
// bram[23628] = 24;
// bram[23629] = 35;
// bram[23630] = 47;
// bram[23631] = 60;
// bram[23632] = 75;
// bram[23633] = 90;
// bram[23634] = 106;
// bram[23635] = 122;
// bram[23636] = 139;
// bram[23637] = 155;
// bram[23638] = 171;
// bram[23639] = 186;
// bram[23640] = 200;
// bram[23641] = 212;
// bram[23642] = 224;
// bram[23643] = 233;
// bram[23644] = 241;
// bram[23645] = 247;
// bram[23646] = 251;
// bram[23647] = 253;
// bram[23648] = 253;
// bram[23649] = 251;
// bram[23650] = 246;
// bram[23651] = 240;
// bram[23652] = 232;
// bram[23653] = 222;
// bram[23654] = 210;
// bram[23655] = 197;
// bram[23656] = 183;
// bram[23657] = 168;
// bram[23658] = 152;
// bram[23659] = 136;
// bram[23660] = 120;
// bram[23661] = 103;
// bram[23662] = 87;
// bram[23663] = 72;
// bram[23664] = 58;
// bram[23665] = 45;
// bram[23666] = 33;
// bram[23667] = 23;
// bram[23668] = 14;
// bram[23669] = 7;
// bram[23670] = 3;
// bram[23671] = 0;
// bram[23672] = 0;
// bram[23673] = 1;
// bram[23674] = 5;
// bram[23675] = 11;
// bram[23676] = 18;
// bram[23677] = 28;
// bram[23678] = 39;
// bram[23679] = 51;
// bram[23680] = 65;
// bram[23681] = 80;
// bram[23682] = 96;
// bram[23683] = 112;
// bram[23684] = 128;
// bram[23685] = 145;
// bram[23686] = 161;
// bram[23687] = 176;
// bram[23688] = 191;
// bram[23689] = 204;
// bram[23690] = 217;
// bram[23691] = 227;
// bram[23692] = 237;
// bram[23693] = 244;
// bram[23694] = 249;
// bram[23695] = 252;
// bram[23696] = 253;
// bram[23697] = 253;
// bram[23698] = 249;
// bram[23699] = 244;
// bram[23700] = 237;
// bram[23701] = 228;
// bram[23702] = 218;
// bram[23703] = 206;
// bram[23704] = 192;
// bram[23705] = 178;
// bram[23706] = 162;
// bram[23707] = 146;
// bram[23708] = 130;
// bram[23709] = 114;
// bram[23710] = 97;
// bram[23711] = 82;
// bram[23712] = 67;
// bram[23713] = 53;
// bram[23714] = 40;
// bram[23715] = 29;
// bram[23716] = 19;
// bram[23717] = 11;
// bram[23718] = 5;
// bram[23719] = 1;
// bram[23720] = 0;
// bram[23721] = 0;
// bram[23722] = 2;
// bram[23723] = 7;
// bram[23724] = 13;
// bram[23725] = 22;
// bram[23726] = 32;
// bram[23727] = 43;
// bram[23728] = 56;
// bram[23729] = 71;
// bram[23730] = 86;
// bram[23731] = 102;
// bram[23732] = 118;
// bram[23733] = 134;
// bram[23734] = 151;
// bram[23735] = 166;
// bram[23736] = 182;
// bram[23737] = 196;
// bram[23738] = 209;
// bram[23739] = 221;
// bram[23740] = 231;
// bram[23741] = 239;
// bram[23742] = 246;
// bram[23743] = 251;
// bram[23744] = 253;
// bram[23745] = 253;
// bram[23746] = 252;
// bram[23747] = 248;
// bram[23748] = 242;
// bram[23749] = 234;
// bram[23750] = 225;
// bram[23751] = 213;
// bram[23752] = 201;
// bram[23753] = 187;
// bram[23754] = 172;
// bram[23755] = 156;
// bram[23756] = 140;
// bram[23757] = 124;
// bram[23758] = 108;
// bram[23759] = 91;
// bram[23760] = 76;
// bram[23761] = 61;
// bram[23762] = 48;
// bram[23763] = 36;
// bram[23764] = 25;
// bram[23765] = 16;
// bram[23766] = 9;
// bram[23767] = 4;
// bram[23768] = 1;
// bram[23769] = 0;
// bram[23770] = 1;
// bram[23771] = 4;
// bram[23772] = 9;
// bram[23773] = 16;
// bram[23774] = 25;
// bram[23775] = 36;
// bram[23776] = 48;
// bram[23777] = 62;
// bram[23778] = 76;
// bram[23779] = 92;
// bram[23780] = 108;
// bram[23781] = 124;
// bram[23782] = 140;
// bram[23783] = 156;
// bram[23784] = 172;
// bram[23785] = 187;
// bram[23786] = 201;
// bram[23787] = 214;
// bram[23788] = 225;
// bram[23789] = 234;
// bram[23790] = 242;
// bram[23791] = 248;
// bram[23792] = 252;
// bram[23793] = 253;
// bram[23794] = 253;
// bram[23795] = 250;
// bram[23796] = 246;
// bram[23797] = 239;
// bram[23798] = 231;
// bram[23799] = 221;
// bram[23800] = 209;
// bram[23801] = 196;
// bram[23802] = 182;
// bram[23803] = 166;
// bram[23804] = 150;
// bram[23805] = 134;
// bram[23806] = 118;
// bram[23807] = 102;
// bram[23808] = 86;
// bram[23809] = 71;
// bram[23810] = 56;
// bram[23811] = 43;
// bram[23812] = 32;
// bram[23813] = 22;
// bram[23814] = 13;
// bram[23815] = 7;
// bram[23816] = 2;
// bram[23817] = 0;
// bram[23818] = 0;
// bram[23819] = 1;
// bram[23820] = 5;
// bram[23821] = 11;
// bram[23822] = 19;
// bram[23823] = 29;
// bram[23824] = 40;
// bram[23825] = 53;
// bram[23826] = 67;
// bram[23827] = 82;
// bram[23828] = 97;
// bram[23829] = 114;
// bram[23830] = 130;
// bram[23831] = 146;
// bram[23832] = 162;
// bram[23833] = 178;
// bram[23834] = 192;
// bram[23835] = 206;
// bram[23836] = 218;
// bram[23837] = 228;
// bram[23838] = 237;
// bram[23839] = 244;
// bram[23840] = 250;
// bram[23841] = 253;
// bram[23842] = 253;
// bram[23843] = 252;
// bram[23844] = 249;
// bram[23845] = 244;
// bram[23846] = 236;
// bram[23847] = 227;
// bram[23848] = 217;
// bram[23849] = 204;
// bram[23850] = 191;
// bram[23851] = 176;
// bram[23852] = 161;
// bram[23853] = 145;
// bram[23854] = 128;
// bram[23855] = 112;
// bram[23856] = 96;
// bram[23857] = 80;
// bram[23858] = 65;
// bram[23859] = 51;
// bram[23860] = 39;
// bram[23861] = 28;
// bram[23862] = 18;
// bram[23863] = 11;
// bram[23864] = 5;
// bram[23865] = 1;
// bram[23866] = 0;
// bram[23867] = 0;
// bram[23868] = 3;
// bram[23869] = 7;
// bram[23870] = 14;
// bram[23871] = 23;
// bram[23872] = 33;
// bram[23873] = 45;
// bram[23874] = 58;
// bram[23875] = 72;
// bram[23876] = 87;
// bram[23877] = 103;
// bram[23878] = 120;
// bram[23879] = 136;
// bram[23880] = 152;
// bram[23881] = 168;
// bram[23882] = 183;
// bram[23883] = 197;
// bram[23884] = 210;
// bram[23885] = 222;
// bram[23886] = 232;
// bram[23887] = 240;
// bram[23888] = 247;
// bram[23889] = 251;
// bram[23890] = 253;
// bram[23891] = 253;
// bram[23892] = 251;
// bram[23893] = 247;
// bram[23894] = 241;
// bram[23895] = 233;
// bram[23896] = 224;
// bram[23897] = 212;
// bram[23898] = 199;
// bram[23899] = 185;
// bram[23900] = 170;
// bram[23901] = 155;
// bram[23902] = 139;
// bram[23903] = 122;
// bram[23904] = 106;
// bram[23905] = 90;
// bram[23906] = 75;
// bram[23907] = 60;
// bram[23908] = 47;
// bram[23909] = 35;
// bram[23910] = 24;
// bram[23911] = 15;
// bram[23912] = 8;
// bram[23913] = 3;
// bram[23914] = 0;
// bram[23915] = 0;
// bram[23916] = 1;
// bram[23917] = 4;
// bram[23918] = 10;
// bram[23919] = 17;
// bram[23920] = 26;
// bram[23921] = 37;
// bram[23922] = 49;
// bram[23923] = 63;
// bram[23924] = 78;
// bram[23925] = 93;
// bram[23926] = 109;
// bram[23927] = 126;
// bram[23928] = 142;
// bram[23929] = 158;
// bram[23930] = 174;
// bram[23931] = 189;
// bram[23932] = 202;
// bram[23933] = 215;
// bram[23934] = 226;
// bram[23935] = 235;
// bram[23936] = 243;
// bram[23937] = 248;
// bram[23938] = 252;
// bram[23939] = 253;
// bram[23940] = 253;
// bram[23941] = 250;
// bram[23942] = 245;
// bram[23943] = 239;
// bram[23944] = 230;
// bram[23945] = 220;
// bram[23946] = 208;
// bram[23947] = 194;
// bram[23948] = 180;
// bram[23949] = 165;
// bram[23950] = 149;
// bram[23951] = 133;
// bram[23952] = 116;
// bram[23953] = 100;
// bram[23954] = 84;
// bram[23955] = 69;
// bram[23956] = 55;
// bram[23957] = 42;
// bram[23958] = 31;
// bram[23959] = 21;
// bram[23960] = 12;
// bram[23961] = 6;
// bram[23962] = 2;
// bram[23963] = 0;
// bram[23964] = 0;
// bram[23965] = 2;
// bram[23966] = 6;
// bram[23967] = 12;
// bram[23968] = 20;
// bram[23969] = 30;
// bram[23970] = 41;
// bram[23971] = 54;
// bram[23972] = 68;
// bram[23973] = 83;
// bram[23974] = 99;
// bram[23975] = 115;
// bram[23976] = 132;
// bram[23977] = 148;
// bram[23978] = 164;
// bram[23979] = 179;
// bram[23980] = 194;
// bram[23981] = 207;
// bram[23982] = 219;
// bram[23983] = 229;
// bram[23984] = 238;
// bram[23985] = 245;
// bram[23986] = 250;
// bram[23987] = 253;
// bram[23988] = 253;
// bram[23989] = 252;
// bram[23990] = 249;
// bram[23991] = 243;
// bram[23992] = 236;
// bram[23993] = 226;
// bram[23994] = 215;
// bram[23995] = 203;
// bram[23996] = 189;
// bram[23997] = 175;
// bram[23998] = 159;
// bram[23999] = 143;
// bram[24000] = 127;
// bram[24001] = 144;
// bram[24002] = 161;
// bram[24003] = 177;
// bram[24004] = 193;
// bram[24005] = 207;
// bram[24006] = 220;
// bram[24007] = 230;
// bram[24008] = 239;
// bram[24009] = 246;
// bram[24010] = 251;
// bram[24011] = 253;
// bram[24012] = 253;
// bram[24013] = 251;
// bram[24014] = 246;
// bram[24015] = 239;
// bram[24016] = 230;
// bram[24017] = 219;
// bram[24018] = 206;
// bram[24019] = 192;
// bram[24020] = 176;
// bram[24021] = 160;
// bram[24022] = 143;
// bram[24023] = 125;
// bram[24024] = 108;
// bram[24025] = 91;
// bram[24026] = 75;
// bram[24027] = 59;
// bram[24028] = 45;
// bram[24029] = 33;
// bram[24030] = 22;
// bram[24031] = 13;
// bram[24032] = 6;
// bram[24033] = 2;
// bram[24034] = 0;
// bram[24035] = 0;
// bram[24036] = 3;
// bram[24037] = 8;
// bram[24038] = 15;
// bram[24039] = 24;
// bram[24040] = 35;
// bram[24041] = 48;
// bram[24042] = 63;
// bram[24043] = 78;
// bram[24044] = 95;
// bram[24045] = 112;
// bram[24046] = 129;
// bram[24047] = 147;
// bram[24048] = 163;
// bram[24049] = 180;
// bram[24050] = 195;
// bram[24051] = 209;
// bram[24052] = 221;
// bram[24053] = 232;
// bram[24054] = 241;
// bram[24055] = 247;
// bram[24056] = 251;
// bram[24057] = 253;
// bram[24058] = 253;
// bram[24059] = 250;
// bram[24060] = 245;
// bram[24061] = 238;
// bram[24062] = 228;
// bram[24063] = 217;
// bram[24064] = 204;
// bram[24065] = 189;
// bram[24066] = 174;
// bram[24067] = 157;
// bram[24068] = 140;
// bram[24069] = 122;
// bram[24070] = 105;
// bram[24071] = 88;
// bram[24072] = 72;
// bram[24073] = 57;
// bram[24074] = 43;
// bram[24075] = 31;
// bram[24076] = 20;
// bram[24077] = 12;
// bram[24078] = 5;
// bram[24079] = 1;
// bram[24080] = 0;
// bram[24081] = 0;
// bram[24082] = 3;
// bram[24083] = 9;
// bram[24084] = 16;
// bram[24085] = 26;
// bram[24086] = 37;
// bram[24087] = 50;
// bram[24088] = 65;
// bram[24089] = 81;
// bram[24090] = 97;
// bram[24091] = 114;
// bram[24092] = 132;
// bram[24093] = 149;
// bram[24094] = 166;
// bram[24095] = 182;
// bram[24096] = 197;
// bram[24097] = 211;
// bram[24098] = 223;
// bram[24099] = 233;
// bram[24100] = 242;
// bram[24101] = 248;
// bram[24102] = 252;
// bram[24103] = 253;
// bram[24104] = 253;
// bram[24105] = 249;
// bram[24106] = 244;
// bram[24107] = 236;
// bram[24108] = 226;
// bram[24109] = 215;
// bram[24110] = 202;
// bram[24111] = 187;
// bram[24112] = 171;
// bram[24113] = 154;
// bram[24114] = 137;
// bram[24115] = 120;
// bram[24116] = 103;
// bram[24117] = 86;
// bram[24118] = 70;
// bram[24119] = 55;
// bram[24120] = 41;
// bram[24121] = 29;
// bram[24122] = 19;
// bram[24123] = 11;
// bram[24124] = 5;
// bram[24125] = 1;
// bram[24126] = 0;
// bram[24127] = 1;
// bram[24128] = 4;
// bram[24129] = 10;
// bram[24130] = 17;
// bram[24131] = 27;
// bram[24132] = 39;
// bram[24133] = 53;
// bram[24134] = 67;
// bram[24135] = 83;
// bram[24136] = 100;
// bram[24137] = 117;
// bram[24138] = 135;
// bram[24139] = 152;
// bram[24140] = 169;
// bram[24141] = 185;
// bram[24142] = 199;
// bram[24143] = 213;
// bram[24144] = 225;
// bram[24145] = 235;
// bram[24146] = 243;
// bram[24147] = 249;
// bram[24148] = 252;
// bram[24149] = 253;
// bram[24150] = 252;
// bram[24151] = 249;
// bram[24152] = 243;
// bram[24153] = 235;
// bram[24154] = 225;
// bram[24155] = 213;
// bram[24156] = 199;
// bram[24157] = 184;
// bram[24158] = 168;
// bram[24159] = 152;
// bram[24160] = 134;
// bram[24161] = 117;
// bram[24162] = 100;
// bram[24163] = 83;
// bram[24164] = 67;
// bram[24165] = 52;
// bram[24166] = 39;
// bram[24167] = 27;
// bram[24168] = 17;
// bram[24169] = 10;
// bram[24170] = 4;
// bram[24171] = 1;
// bram[24172] = 0;
// bram[24173] = 1;
// bram[24174] = 5;
// bram[24175] = 11;
// bram[24176] = 19;
// bram[24177] = 29;
// bram[24178] = 41;
// bram[24179] = 55;
// bram[24180] = 70;
// bram[24181] = 86;
// bram[24182] = 103;
// bram[24183] = 120;
// bram[24184] = 137;
// bram[24185] = 154;
// bram[24186] = 171;
// bram[24187] = 187;
// bram[24188] = 202;
// bram[24189] = 215;
// bram[24190] = 227;
// bram[24191] = 236;
// bram[24192] = 244;
// bram[24193] = 249;
// bram[24194] = 253;
// bram[24195] = 253;
// bram[24196] = 252;
// bram[24197] = 248;
// bram[24198] = 242;
// bram[24199] = 233;
// bram[24200] = 223;
// bram[24201] = 211;
// bram[24202] = 197;
// bram[24203] = 182;
// bram[24204] = 166;
// bram[24205] = 149;
// bram[24206] = 132;
// bram[24207] = 114;
// bram[24208] = 97;
// bram[24209] = 81;
// bram[24210] = 65;
// bram[24211] = 50;
// bram[24212] = 37;
// bram[24213] = 26;
// bram[24214] = 16;
// bram[24215] = 9;
// bram[24216] = 3;
// bram[24217] = 0;
// bram[24218] = 0;
// bram[24219] = 1;
// bram[24220] = 5;
// bram[24221] = 12;
// bram[24222] = 20;
// bram[24223] = 31;
// bram[24224] = 43;
// bram[24225] = 57;
// bram[24226] = 72;
// bram[24227] = 88;
// bram[24228] = 105;
// bram[24229] = 123;
// bram[24230] = 140;
// bram[24231] = 157;
// bram[24232] = 174;
// bram[24233] = 189;
// bram[24234] = 204;
// bram[24235] = 217;
// bram[24236] = 228;
// bram[24237] = 238;
// bram[24238] = 245;
// bram[24239] = 250;
// bram[24240] = 253;
// bram[24241] = 253;
// bram[24242] = 251;
// bram[24243] = 247;
// bram[24244] = 241;
// bram[24245] = 232;
// bram[24246] = 221;
// bram[24247] = 209;
// bram[24248] = 195;
// bram[24249] = 180;
// bram[24250] = 163;
// bram[24251] = 146;
// bram[24252] = 129;
// bram[24253] = 112;
// bram[24254] = 95;
// bram[24255] = 78;
// bram[24256] = 63;
// bram[24257] = 48;
// bram[24258] = 35;
// bram[24259] = 24;
// bram[24260] = 15;
// bram[24261] = 8;
// bram[24262] = 3;
// bram[24263] = 0;
// bram[24264] = 0;
// bram[24265] = 2;
// bram[24266] = 6;
// bram[24267] = 13;
// bram[24268] = 22;
// bram[24269] = 33;
// bram[24270] = 45;
// bram[24271] = 59;
// bram[24272] = 75;
// bram[24273] = 91;
// bram[24274] = 108;
// bram[24275] = 125;
// bram[24276] = 143;
// bram[24277] = 160;
// bram[24278] = 176;
// bram[24279] = 192;
// bram[24280] = 206;
// bram[24281] = 219;
// bram[24282] = 230;
// bram[24283] = 239;
// bram[24284] = 246;
// bram[24285] = 251;
// bram[24286] = 253;
// bram[24287] = 253;
// bram[24288] = 251;
// bram[24289] = 246;
// bram[24290] = 239;
// bram[24291] = 230;
// bram[24292] = 219;
// bram[24293] = 207;
// bram[24294] = 193;
// bram[24295] = 177;
// bram[24296] = 161;
// bram[24297] = 144;
// bram[24298] = 126;
// bram[24299] = 109;
// bram[24300] = 92;
// bram[24301] = 76;
// bram[24302] = 60;
// bram[24303] = 46;
// bram[24304] = 33;
// bram[24305] = 22;
// bram[24306] = 13;
// bram[24307] = 7;
// bram[24308] = 2;
// bram[24309] = 0;
// bram[24310] = 0;
// bram[24311] = 2;
// bram[24312] = 7;
// bram[24313] = 14;
// bram[24314] = 23;
// bram[24315] = 34;
// bram[24316] = 47;
// bram[24317] = 62;
// bram[24318] = 77;
// bram[24319] = 94;
// bram[24320] = 111;
// bram[24321] = 128;
// bram[24322] = 145;
// bram[24323] = 162;
// bram[24324] = 179;
// bram[24325] = 194;
// bram[24326] = 208;
// bram[24327] = 221;
// bram[24328] = 231;
// bram[24329] = 240;
// bram[24330] = 247;
// bram[24331] = 251;
// bram[24332] = 253;
// bram[24333] = 253;
// bram[24334] = 250;
// bram[24335] = 245;
// bram[24336] = 238;
// bram[24337] = 229;
// bram[24338] = 218;
// bram[24339] = 205;
// bram[24340] = 190;
// bram[24341] = 175;
// bram[24342] = 158;
// bram[24343] = 141;
// bram[24344] = 124;
// bram[24345] = 106;
// bram[24346] = 89;
// bram[24347] = 73;
// bram[24348] = 58;
// bram[24349] = 44;
// bram[24350] = 32;
// bram[24351] = 21;
// bram[24352] = 12;
// bram[24353] = 6;
// bram[24354] = 2;
// bram[24355] = 0;
// bram[24356] = 0;
// bram[24357] = 3;
// bram[24358] = 8;
// bram[24359] = 15;
// bram[24360] = 25;
// bram[24361] = 36;
// bram[24362] = 49;
// bram[24363] = 64;
// bram[24364] = 80;
// bram[24365] = 96;
// bram[24366] = 113;
// bram[24367] = 131;
// bram[24368] = 148;
// bram[24369] = 165;
// bram[24370] = 181;
// bram[24371] = 196;
// bram[24372] = 210;
// bram[24373] = 222;
// bram[24374] = 233;
// bram[24375] = 241;
// bram[24376] = 248;
// bram[24377] = 252;
// bram[24378] = 253;
// bram[24379] = 253;
// bram[24380] = 250;
// bram[24381] = 244;
// bram[24382] = 237;
// bram[24383] = 227;
// bram[24384] = 216;
// bram[24385] = 203;
// bram[24386] = 188;
// bram[24387] = 172;
// bram[24388] = 156;
// bram[24389] = 138;
// bram[24390] = 121;
// bram[24391] = 104;
// bram[24392] = 87;
// bram[24393] = 71;
// bram[24394] = 56;
// bram[24395] = 42;
// bram[24396] = 30;
// bram[24397] = 19;
// bram[24398] = 11;
// bram[24399] = 5;
// bram[24400] = 1;
// bram[24401] = 0;
// bram[24402] = 0;
// bram[24403] = 4;
// bram[24404] = 9;
// bram[24405] = 17;
// bram[24406] = 27;
// bram[24407] = 38;
// bram[24408] = 52;
// bram[24409] = 66;
// bram[24410] = 82;
// bram[24411] = 99;
// bram[24412] = 116;
// bram[24413] = 133;
// bram[24414] = 151;
// bram[24415] = 167;
// bram[24416] = 183;
// bram[24417] = 198;
// bram[24418] = 212;
// bram[24419] = 224;
// bram[24420] = 234;
// bram[24421] = 242;
// bram[24422] = 248;
// bram[24423] = 252;
// bram[24424] = 253;
// bram[24425] = 252;
// bram[24426] = 249;
// bram[24427] = 243;
// bram[24428] = 236;
// bram[24429] = 226;
// bram[24430] = 214;
// bram[24431] = 200;
// bram[24432] = 186;
// bram[24433] = 170;
// bram[24434] = 153;
// bram[24435] = 136;
// bram[24436] = 118;
// bram[24437] = 101;
// bram[24438] = 84;
// bram[24439] = 68;
// bram[24440] = 53;
// bram[24441] = 40;
// bram[24442] = 28;
// bram[24443] = 18;
// bram[24444] = 10;
// bram[24445] = 4;
// bram[24446] = 1;
// bram[24447] = 0;
// bram[24448] = 1;
// bram[24449] = 4;
// bram[24450] = 10;
// bram[24451] = 18;
// bram[24452] = 28;
// bram[24453] = 40;
// bram[24454] = 54;
// bram[24455] = 69;
// bram[24456] = 85;
// bram[24457] = 101;
// bram[24458] = 119;
// bram[24459] = 136;
// bram[24460] = 153;
// bram[24461] = 170;
// bram[24462] = 186;
// bram[24463] = 201;
// bram[24464] = 214;
// bram[24465] = 226;
// bram[24466] = 236;
// bram[24467] = 244;
// bram[24468] = 249;
// bram[24469] = 253;
// bram[24470] = 253;
// bram[24471] = 252;
// bram[24472] = 248;
// bram[24473] = 242;
// bram[24474] = 234;
// bram[24475] = 224;
// bram[24476] = 212;
// bram[24477] = 198;
// bram[24478] = 183;
// bram[24479] = 167;
// bram[24480] = 150;
// bram[24481] = 133;
// bram[24482] = 116;
// bram[24483] = 98;
// bram[24484] = 82;
// bram[24485] = 66;
// bram[24486] = 51;
// bram[24487] = 38;
// bram[24488] = 26;
// bram[24489] = 17;
// bram[24490] = 9;
// bram[24491] = 4;
// bram[24492] = 0;
// bram[24493] = 0;
// bram[24494] = 1;
// bram[24495] = 5;
// bram[24496] = 11;
// bram[24497] = 20;
// bram[24498] = 30;
// bram[24499] = 42;
// bram[24500] = 56;
// bram[24501] = 71;
// bram[24502] = 87;
// bram[24503] = 104;
// bram[24504] = 121;
// bram[24505] = 139;
// bram[24506] = 156;
// bram[24507] = 172;
// bram[24508] = 188;
// bram[24509] = 203;
// bram[24510] = 216;
// bram[24511] = 227;
// bram[24512] = 237;
// bram[24513] = 245;
// bram[24514] = 250;
// bram[24515] = 253;
// bram[24516] = 253;
// bram[24517] = 252;
// bram[24518] = 248;
// bram[24519] = 241;
// bram[24520] = 233;
// bram[24521] = 222;
// bram[24522] = 210;
// bram[24523] = 196;
// bram[24524] = 181;
// bram[24525] = 165;
// bram[24526] = 148;
// bram[24527] = 130;
// bram[24528] = 113;
// bram[24529] = 96;
// bram[24530] = 79;
// bram[24531] = 64;
// bram[24532] = 49;
// bram[24533] = 36;
// bram[24534] = 25;
// bram[24535] = 15;
// bram[24536] = 8;
// bram[24537] = 3;
// bram[24538] = 0;
// bram[24539] = 0;
// bram[24540] = 2;
// bram[24541] = 6;
// bram[24542] = 12;
// bram[24543] = 21;
// bram[24544] = 32;
// bram[24545] = 44;
// bram[24546] = 58;
// bram[24547] = 73;
// bram[24548] = 90;
// bram[24549] = 107;
// bram[24550] = 124;
// bram[24551] = 141;
// bram[24552] = 158;
// bram[24553] = 175;
// bram[24554] = 191;
// bram[24555] = 205;
// bram[24556] = 218;
// bram[24557] = 229;
// bram[24558] = 238;
// bram[24559] = 245;
// bram[24560] = 250;
// bram[24561] = 253;
// bram[24562] = 253;
// bram[24563] = 251;
// bram[24564] = 247;
// bram[24565] = 240;
// bram[24566] = 231;
// bram[24567] = 220;
// bram[24568] = 208;
// bram[24569] = 194;
// bram[24570] = 178;
// bram[24571] = 162;
// bram[24572] = 145;
// bram[24573] = 128;
// bram[24574] = 110;
// bram[24575] = 93;
// bram[24576] = 77;
// bram[24577] = 61;
// bram[24578] = 47;
// bram[24579] = 34;
// bram[24580] = 23;
// bram[24581] = 14;
// bram[24582] = 7;
// bram[24583] = 2;
// bram[24584] = 0;
// bram[24585] = 0;
// bram[24586] = 2;
// bram[24587] = 7;
// bram[24588] = 14;
// bram[24589] = 23;
// bram[24590] = 34;
// bram[24591] = 46;
// bram[24592] = 60;
// bram[24593] = 76;
// bram[24594] = 92;
// bram[24595] = 109;
// bram[24596] = 127;
// bram[24597] = 144;
// bram[24598] = 161;
// bram[24599] = 177;
// bram[24600] = 193;
// bram[24601] = 207;
// bram[24602] = 220;
// bram[24603] = 231;
// bram[24604] = 240;
// bram[24605] = 246;
// bram[24606] = 251;
// bram[24607] = 253;
// bram[24608] = 253;
// bram[24609] = 251;
// bram[24610] = 246;
// bram[24611] = 239;
// bram[24612] = 230;
// bram[24613] = 218;
// bram[24614] = 206;
// bram[24615] = 191;
// bram[24616] = 176;
// bram[24617] = 159;
// bram[24618] = 142;
// bram[24619] = 125;
// bram[24620] = 108;
// bram[24621] = 91;
// bram[24622] = 74;
// bram[24623] = 59;
// bram[24624] = 45;
// bram[24625] = 32;
// bram[24626] = 22;
// bram[24627] = 13;
// bram[24628] = 6;
// bram[24629] = 2;
// bram[24630] = 0;
// bram[24631] = 0;
// bram[24632] = 3;
// bram[24633] = 8;
// bram[24634] = 15;
// bram[24635] = 24;
// bram[24636] = 35;
// bram[24637] = 48;
// bram[24638] = 63;
// bram[24639] = 78;
// bram[24640] = 95;
// bram[24641] = 112;
// bram[24642] = 129;
// bram[24643] = 147;
// bram[24644] = 164;
// bram[24645] = 180;
// bram[24646] = 195;
// bram[24647] = 209;
// bram[24648] = 221;
// bram[24649] = 232;
// bram[24650] = 241;
// bram[24651] = 247;
// bram[24652] = 252;
// bram[24653] = 253;
// bram[24654] = 253;
// bram[24655] = 250;
// bram[24656] = 245;
// bram[24657] = 237;
// bram[24658] = 228;
// bram[24659] = 217;
// bram[24660] = 204;
// bram[24661] = 189;
// bram[24662] = 173;
// bram[24663] = 157;
// bram[24664] = 140;
// bram[24665] = 122;
// bram[24666] = 105;
// bram[24667] = 88;
// bram[24668] = 72;
// bram[24669] = 57;
// bram[24670] = 43;
// bram[24671] = 31;
// bram[24672] = 20;
// bram[24673] = 12;
// bram[24674] = 5;
// bram[24675] = 1;
// bram[24676] = 0;
// bram[24677] = 0;
// bram[24678] = 3;
// bram[24679] = 9;
// bram[24680] = 16;
// bram[24681] = 26;
// bram[24682] = 37;
// bram[24683] = 51;
// bram[24684] = 65;
// bram[24685] = 81;
// bram[24686] = 98;
// bram[24687] = 115;
// bram[24688] = 132;
// bram[24689] = 149;
// bram[24690] = 166;
// bram[24691] = 182;
// bram[24692] = 197;
// bram[24693] = 211;
// bram[24694] = 223;
// bram[24695] = 234;
// bram[24696] = 242;
// bram[24697] = 248;
// bram[24698] = 252;
// bram[24699] = 253;
// bram[24700] = 253;
// bram[24701] = 249;
// bram[24702] = 244;
// bram[24703] = 236;
// bram[24704] = 226;
// bram[24705] = 215;
// bram[24706] = 201;
// bram[24707] = 187;
// bram[24708] = 171;
// bram[24709] = 154;
// bram[24710] = 137;
// bram[24711] = 120;
// bram[24712] = 102;
// bram[24713] = 86;
// bram[24714] = 69;
// bram[24715] = 54;
// bram[24716] = 41;
// bram[24717] = 29;
// bram[24718] = 19;
// bram[24719] = 11;
// bram[24720] = 5;
// bram[24721] = 1;
// bram[24722] = 0;
// bram[24723] = 1;
// bram[24724] = 4;
// bram[24725] = 10;
// bram[24726] = 18;
// bram[24727] = 27;
// bram[24728] = 39;
// bram[24729] = 53;
// bram[24730] = 68;
// bram[24731] = 83;
// bram[24732] = 100;
// bram[24733] = 117;
// bram[24734] = 135;
// bram[24735] = 152;
// bram[24736] = 169;
// bram[24737] = 185;
// bram[24738] = 200;
// bram[24739] = 213;
// bram[24740] = 225;
// bram[24741] = 235;
// bram[24742] = 243;
// bram[24743] = 249;
// bram[24744] = 252;
// bram[24745] = 253;
// bram[24746] = 252;
// bram[24747] = 249;
// bram[24748] = 243;
// bram[24749] = 235;
// bram[24750] = 225;
// bram[24751] = 213;
// bram[24752] = 199;
// bram[24753] = 184;
// bram[24754] = 168;
// bram[24755] = 152;
// bram[24756] = 134;
// bram[24757] = 117;
// bram[24758] = 100;
// bram[24759] = 83;
// bram[24760] = 67;
// bram[24761] = 52;
// bram[24762] = 39;
// bram[24763] = 27;
// bram[24764] = 17;
// bram[24765] = 9;
// bram[24766] = 4;
// bram[24767] = 0;
// bram[24768] = 0;
// bram[24769] = 1;
// bram[24770] = 5;
// bram[24771] = 11;
// bram[24772] = 19;
// bram[24773] = 29;
// bram[24774] = 41;
// bram[24775] = 55;
// bram[24776] = 70;
// bram[24777] = 86;
// bram[24778] = 103;
// bram[24779] = 120;
// bram[24780] = 137;
// bram[24781] = 155;
// bram[24782] = 171;
// bram[24783] = 187;
// bram[24784] = 202;
// bram[24785] = 215;
// bram[24786] = 227;
// bram[24787] = 236;
// bram[24788] = 244;
// bram[24789] = 250;
// bram[24790] = 253;
// bram[24791] = 253;
// bram[24792] = 252;
// bram[24793] = 248;
// bram[24794] = 242;
// bram[24795] = 233;
// bram[24796] = 223;
// bram[24797] = 211;
// bram[24798] = 197;
// bram[24799] = 182;
// bram[24800] = 166;
// bram[24801] = 149;
// bram[24802] = 132;
// bram[24803] = 114;
// bram[24804] = 97;
// bram[24805] = 80;
// bram[24806] = 65;
// bram[24807] = 50;
// bram[24808] = 37;
// bram[24809] = 26;
// bram[24810] = 16;
// bram[24811] = 8;
// bram[24812] = 3;
// bram[24813] = 0;
// bram[24814] = 0;
// bram[24815] = 1;
// bram[24816] = 5;
// bram[24817] = 12;
// bram[24818] = 20;
// bram[24819] = 31;
// bram[24820] = 43;
// bram[24821] = 57;
// bram[24822] = 72;
// bram[24823] = 89;
// bram[24824] = 105;
// bram[24825] = 123;
// bram[24826] = 140;
// bram[24827] = 157;
// bram[24828] = 174;
// bram[24829] = 189;
// bram[24830] = 204;
// bram[24831] = 217;
// bram[24832] = 228;
// bram[24833] = 238;
// bram[24834] = 245;
// bram[24835] = 250;
// bram[24836] = 253;
// bram[24837] = 253;
// bram[24838] = 251;
// bram[24839] = 247;
// bram[24840] = 241;
// bram[24841] = 232;
// bram[24842] = 221;
// bram[24843] = 209;
// bram[24844] = 195;
// bram[24845] = 179;
// bram[24846] = 163;
// bram[24847] = 146;
// bram[24848] = 129;
// bram[24849] = 112;
// bram[24850] = 94;
// bram[24851] = 78;
// bram[24852] = 62;
// bram[24853] = 48;
// bram[24854] = 35;
// bram[24855] = 24;
// bram[24856] = 15;
// bram[24857] = 7;
// bram[24858] = 3;
// bram[24859] = 0;
// bram[24860] = 0;
// bram[24861] = 2;
// bram[24862] = 6;
// bram[24863] = 13;
// bram[24864] = 22;
// bram[24865] = 33;
// bram[24866] = 45;
// bram[24867] = 59;
// bram[24868] = 75;
// bram[24869] = 91;
// bram[24870] = 108;
// bram[24871] = 125;
// bram[24872] = 143;
// bram[24873] = 160;
// bram[24874] = 176;
// bram[24875] = 192;
// bram[24876] = 206;
// bram[24877] = 219;
// bram[24878] = 230;
// bram[24879] = 239;
// bram[24880] = 246;
// bram[24881] = 251;
// bram[24882] = 253;
// bram[24883] = 253;
// bram[24884] = 251;
// bram[24885] = 246;
// bram[24886] = 239;
// bram[24887] = 230;
// bram[24888] = 219;
// bram[24889] = 207;
// bram[24890] = 192;
// bram[24891] = 177;
// bram[24892] = 161;
// bram[24893] = 144;
// bram[24894] = 126;
// bram[24895] = 109;
// bram[24896] = 92;
// bram[24897] = 75;
// bram[24898] = 60;
// bram[24899] = 46;
// bram[24900] = 33;
// bram[24901] = 22;
// bram[24902] = 13;
// bram[24903] = 7;
// bram[24904] = 2;
// bram[24905] = 0;
// bram[24906] = 0;
// bram[24907] = 2;
// bram[24908] = 7;
// bram[24909] = 14;
// bram[24910] = 23;
// bram[24911] = 35;
// bram[24912] = 47;
// bram[24913] = 62;
// bram[24914] = 77;
// bram[24915] = 94;
// bram[24916] = 111;
// bram[24917] = 128;
// bram[24918] = 145;
// bram[24919] = 162;
// bram[24920] = 179;
// bram[24921] = 194;
// bram[24922] = 208;
// bram[24923] = 221;
// bram[24924] = 231;
// bram[24925] = 240;
// bram[24926] = 247;
// bram[24927] = 251;
// bram[24928] = 253;
// bram[24929] = 253;
// bram[24930] = 250;
// bram[24931] = 245;
// bram[24932] = 238;
// bram[24933] = 229;
// bram[24934] = 217;
// bram[24935] = 205;
// bram[24936] = 190;
// bram[24937] = 175;
// bram[24938] = 158;
// bram[24939] = 141;
// bram[24940] = 124;
// bram[24941] = 106;
// bram[24942] = 89;
// bram[24943] = 73;
// bram[24944] = 58;
// bram[24945] = 44;
// bram[24946] = 31;
// bram[24947] = 21;
// bram[24948] = 12;
// bram[24949] = 6;
// bram[24950] = 1;
// bram[24951] = 0;
// bram[24952] = 0;
// bram[24953] = 3;
// bram[24954] = 8;
// bram[24955] = 16;
// bram[24956] = 25;
// bram[24957] = 36;
// bram[24958] = 50;
// bram[24959] = 64;
// bram[24960] = 80;
// bram[24961] = 96;
// bram[24962] = 113;
// bram[24963] = 131;
// bram[24964] = 148;
// bram[24965] = 165;
// bram[24966] = 181;
// bram[24967] = 196;
// bram[24968] = 210;
// bram[24969] = 222;
// bram[24970] = 233;
// bram[24971] = 241;
// bram[24972] = 248;
// bram[24973] = 252;
// bram[24974] = 253;
// bram[24975] = 253;
// bram[24976] = 250;
// bram[24977] = 244;
// bram[24978] = 237;
// bram[24979] = 227;
// bram[24980] = 216;
// bram[24981] = 202;
// bram[24982] = 188;
// bram[24983] = 172;
// bram[24984] = 155;
// bram[24985] = 138;
// bram[24986] = 121;
// bram[24987] = 104;
// bram[24988] = 87;
// bram[24989] = 71;
// bram[24990] = 56;
// bram[24991] = 42;
// bram[24992] = 30;
// bram[24993] = 19;
// bram[24994] = 11;
// bram[24995] = 5;
// bram[24996] = 1;
// bram[24997] = 0;
// bram[24998] = 0;
// bram[24999] = 4;
// bram[25000] = 9;
// bram[25001] = 17;
// bram[25002] = 27;
// bram[25003] = 38;
// bram[25004] = 52;
// bram[25005] = 66;
// bram[25006] = 82;
// bram[25007] = 99;
// bram[25008] = 116;
// bram[25009] = 134;
// bram[25010] = 151;
// bram[25011] = 168;
// bram[25012] = 184;
// bram[25013] = 199;
// bram[25014] = 212;
// bram[25015] = 224;
// bram[25016] = 234;
// bram[25017] = 243;
// bram[25018] = 248;
// bram[25019] = 252;
// bram[25020] = 253;
// bram[25021] = 252;
// bram[25022] = 249;
// bram[25023] = 243;
// bram[25024] = 235;
// bram[25025] = 225;
// bram[25026] = 214;
// bram[25027] = 200;
// bram[25028] = 185;
// bram[25029] = 169;
// bram[25030] = 153;
// bram[25031] = 136;
// bram[25032] = 118;
// bram[25033] = 101;
// bram[25034] = 84;
// bram[25035] = 68;
// bram[25036] = 53;
// bram[25037] = 40;
// bram[25038] = 28;
// bram[25039] = 18;
// bram[25040] = 10;
// bram[25041] = 4;
// bram[25042] = 1;
// bram[25043] = 0;
// bram[25044] = 1;
// bram[25045] = 4;
// bram[25046] = 10;
// bram[25047] = 18;
// bram[25048] = 28;
// bram[25049] = 40;
// bram[25050] = 54;
// bram[25051] = 69;
// bram[25052] = 85;
// bram[25053] = 102;
// bram[25054] = 119;
// bram[25055] = 136;
// bram[25056] = 153;
// bram[25057] = 170;
// bram[25058] = 186;
// bram[25059] = 201;
// bram[25060] = 214;
// bram[25061] = 226;
// bram[25062] = 236;
// bram[25063] = 244;
// bram[25064] = 249;
// bram[25065] = 253;
// bram[25066] = 253;
// bram[25067] = 252;
// bram[25068] = 248;
// bram[25069] = 242;
// bram[25070] = 234;
// bram[25071] = 224;
// bram[25072] = 212;
// bram[25073] = 198;
// bram[25074] = 183;
// bram[25075] = 167;
// bram[25076] = 150;
// bram[25077] = 133;
// bram[25078] = 115;
// bram[25079] = 98;
// bram[25080] = 82;
// bram[25081] = 66;
// bram[25082] = 51;
// bram[25083] = 38;
// bram[25084] = 26;
// bram[25085] = 17;
// bram[25086] = 9;
// bram[25087] = 3;
// bram[25088] = 0;
// bram[25089] = 0;
// bram[25090] = 1;
// bram[25091] = 5;
// bram[25092] = 11;
// bram[25093] = 20;
// bram[25094] = 30;
// bram[25095] = 42;
// bram[25096] = 56;
// bram[25097] = 71;
// bram[25098] = 87;
// bram[25099] = 104;
// bram[25100] = 122;
// bram[25101] = 139;
// bram[25102] = 156;
// bram[25103] = 173;
// bram[25104] = 188;
// bram[25105] = 203;
// bram[25106] = 216;
// bram[25107] = 228;
// bram[25108] = 237;
// bram[25109] = 245;
// bram[25110] = 250;
// bram[25111] = 253;
// bram[25112] = 253;
// bram[25113] = 252;
// bram[25114] = 247;
// bram[25115] = 241;
// bram[25116] = 233;
// bram[25117] = 222;
// bram[25118] = 210;
// bram[25119] = 196;
// bram[25120] = 181;
// bram[25121] = 164;
// bram[25122] = 147;
// bram[25123] = 130;
// bram[25124] = 113;
// bram[25125] = 96;
// bram[25126] = 79;
// bram[25127] = 63;
// bram[25128] = 49;
// bram[25129] = 36;
// bram[25130] = 25;
// bram[25131] = 15;
// bram[25132] = 8;
// bram[25133] = 3;
// bram[25134] = 0;
// bram[25135] = 0;
// bram[25136] = 2;
// bram[25137] = 6;
// bram[25138] = 12;
// bram[25139] = 21;
// bram[25140] = 32;
// bram[25141] = 44;
// bram[25142] = 58;
// bram[25143] = 74;
// bram[25144] = 90;
// bram[25145] = 107;
// bram[25146] = 124;
// bram[25147] = 142;
// bram[25148] = 159;
// bram[25149] = 175;
// bram[25150] = 191;
// bram[25151] = 205;
// bram[25152] = 218;
// bram[25153] = 229;
// bram[25154] = 238;
// bram[25155] = 246;
// bram[25156] = 250;
// bram[25157] = 253;
// bram[25158] = 253;
// bram[25159] = 251;
// bram[25160] = 247;
// bram[25161] = 240;
// bram[25162] = 231;
// bram[25163] = 220;
// bram[25164] = 208;
// bram[25165] = 193;
// bram[25166] = 178;
// bram[25167] = 162;
// bram[25168] = 145;
// bram[25169] = 127;
// bram[25170] = 110;
// bram[25171] = 93;
// bram[25172] = 77;
// bram[25173] = 61;
// bram[25174] = 47;
// bram[25175] = 34;
// bram[25176] = 23;
// bram[25177] = 14;
// bram[25178] = 7;
// bram[25179] = 2;
// bram[25180] = 0;
// bram[25181] = 0;
// bram[25182] = 2;
// bram[25183] = 7;
// bram[25184] = 14;
// bram[25185] = 23;
// bram[25186] = 34;
// bram[25187] = 46;
// bram[25188] = 61;
// bram[25189] = 76;
// bram[25190] = 93;
// bram[25191] = 110;
// bram[25192] = 127;
// bram[25193] = 144;
// bram[25194] = 161;
// bram[25195] = 178;
// bram[25196] = 193;
// bram[25197] = 207;
// bram[25198] = 220;
// bram[25199] = 231;
// bram[25200] = 240;
// bram[25201] = 246;
// bram[25202] = 251;
// bram[25203] = 253;
// bram[25204] = 253;
// bram[25205] = 251;
// bram[25206] = 246;
// bram[25207] = 239;
// bram[25208] = 229;
// bram[25209] = 218;
// bram[25210] = 206;
// bram[25211] = 191;
// bram[25212] = 176;
// bram[25213] = 159;
// bram[25214] = 142;
// bram[25215] = 125;
// bram[25216] = 107;
// bram[25217] = 90;
// bram[25218] = 74;
// bram[25219] = 59;
// bram[25220] = 45;
// bram[25221] = 32;
// bram[25222] = 22;
// bram[25223] = 13;
// bram[25224] = 6;
// bram[25225] = 2;
// bram[25226] = 0;
// bram[25227] = 0;
// bram[25228] = 3;
// bram[25229] = 8;
// bram[25230] = 15;
// bram[25231] = 24;
// bram[25232] = 36;
// bram[25233] = 49;
// bram[25234] = 63;
// bram[25235] = 79;
// bram[25236] = 95;
// bram[25237] = 112;
// bram[25238] = 130;
// bram[25239] = 147;
// bram[25240] = 164;
// bram[25241] = 180;
// bram[25242] = 195;
// bram[25243] = 209;
// bram[25244] = 222;
// bram[25245] = 232;
// bram[25246] = 241;
// bram[25247] = 247;
// bram[25248] = 252;
// bram[25249] = 253;
// bram[25250] = 253;
// bram[25251] = 250;
// bram[25252] = 245;
// bram[25253] = 237;
// bram[25254] = 228;
// bram[25255] = 216;
// bram[25256] = 203;
// bram[25257] = 189;
// bram[25258] = 173;
// bram[25259] = 157;
// bram[25260] = 139;
// bram[25261] = 122;
// bram[25262] = 105;
// bram[25263] = 88;
// bram[25264] = 72;
// bram[25265] = 57;
// bram[25266] = 43;
// bram[25267] = 30;
// bram[25268] = 20;
// bram[25269] = 12;
// bram[25270] = 5;
// bram[25271] = 1;
// bram[25272] = 0;
// bram[25273] = 0;
// bram[25274] = 3;
// bram[25275] = 9;
// bram[25276] = 16;
// bram[25277] = 26;
// bram[25278] = 37;
// bram[25279] = 51;
// bram[25280] = 65;
// bram[25281] = 81;
// bram[25282] = 98;
// bram[25283] = 115;
// bram[25284] = 132;
// bram[25285] = 150;
// bram[25286] = 166;
// bram[25287] = 183;
// bram[25288] = 198;
// bram[25289] = 211;
// bram[25290] = 223;
// bram[25291] = 234;
// bram[25292] = 242;
// bram[25293] = 248;
// bram[25294] = 252;
// bram[25295] = 253;
// bram[25296] = 253;
// bram[25297] = 249;
// bram[25298] = 244;
// bram[25299] = 236;
// bram[25300] = 226;
// bram[25301] = 215;
// bram[25302] = 201;
// bram[25303] = 186;
// bram[25304] = 171;
// bram[25305] = 154;
// bram[25306] = 137;
// bram[25307] = 119;
// bram[25308] = 102;
// bram[25309] = 85;
// bram[25310] = 69;
// bram[25311] = 54;
// bram[25312] = 41;
// bram[25313] = 29;
// bram[25314] = 19;
// bram[25315] = 10;
// bram[25316] = 4;
// bram[25317] = 1;
// bram[25318] = 0;
// bram[25319] = 1;
// bram[25320] = 4;
// bram[25321] = 10;
// bram[25322] = 18;
// bram[25323] = 28;
// bram[25324] = 39;
// bram[25325] = 53;
// bram[25326] = 68;
// bram[25327] = 84;
// bram[25328] = 100;
// bram[25329] = 118;
// bram[25330] = 135;
// bram[25331] = 152;
// bram[25332] = 169;
// bram[25333] = 185;
// bram[25334] = 200;
// bram[25335] = 213;
// bram[25336] = 225;
// bram[25337] = 235;
// bram[25338] = 243;
// bram[25339] = 249;
// bram[25340] = 252;
// bram[25341] = 253;
// bram[25342] = 252;
// bram[25343] = 249;
// bram[25344] = 243;
// bram[25345] = 235;
// bram[25346] = 225;
// bram[25347] = 213;
// bram[25348] = 199;
// bram[25349] = 184;
// bram[25350] = 168;
// bram[25351] = 151;
// bram[25352] = 134;
// bram[25353] = 117;
// bram[25354] = 99;
// bram[25355] = 83;
// bram[25356] = 67;
// bram[25357] = 52;
// bram[25358] = 39;
// bram[25359] = 27;
// bram[25360] = 17;
// bram[25361] = 9;
// bram[25362] = 4;
// bram[25363] = 0;
// bram[25364] = 0;
// bram[25365] = 1;
// bram[25366] = 5;
// bram[25367] = 11;
// bram[25368] = 19;
// bram[25369] = 29;
// bram[25370] = 41;
// bram[25371] = 55;
// bram[25372] = 70;
// bram[25373] = 86;
// bram[25374] = 103;
// bram[25375] = 120;
// bram[25376] = 138;
// bram[25377] = 155;
// bram[25378] = 171;
// bram[25379] = 187;
// bram[25380] = 202;
// bram[25381] = 215;
// bram[25382] = 227;
// bram[25383] = 236;
// bram[25384] = 244;
// bram[25385] = 250;
// bram[25386] = 253;
// bram[25387] = 253;
// bram[25388] = 252;
// bram[25389] = 248;
// bram[25390] = 242;
// bram[25391] = 233;
// bram[25392] = 223;
// bram[25393] = 211;
// bram[25394] = 197;
// bram[25395] = 182;
// bram[25396] = 166;
// bram[25397] = 149;
// bram[25398] = 131;
// bram[25399] = 114;
// bram[25400] = 97;
// bram[25401] = 80;
// bram[25402] = 65;
// bram[25403] = 50;
// bram[25404] = 37;
// bram[25405] = 25;
// bram[25406] = 16;
// bram[25407] = 8;
// bram[25408] = 3;
// bram[25409] = 0;
// bram[25410] = 0;
// bram[25411] = 1;
// bram[25412] = 6;
// bram[25413] = 12;
// bram[25414] = 21;
// bram[25415] = 31;
// bram[25416] = 43;
// bram[25417] = 57;
// bram[25418] = 73;
// bram[25419] = 89;
// bram[25420] = 106;
// bram[25421] = 123;
// bram[25422] = 140;
// bram[25423] = 157;
// bram[25424] = 174;
// bram[25425] = 190;
// bram[25426] = 204;
// bram[25427] = 217;
// bram[25428] = 228;
// bram[25429] = 238;
// bram[25430] = 245;
// bram[25431] = 250;
// bram[25432] = 253;
// bram[25433] = 253;
// bram[25434] = 251;
// bram[25435] = 247;
// bram[25436] = 240;
// bram[25437] = 232;
// bram[25438] = 221;
// bram[25439] = 209;
// bram[25440] = 195;
// bram[25441] = 179;
// bram[25442] = 163;
// bram[25443] = 146;
// bram[25444] = 129;
// bram[25445] = 111;
// bram[25446] = 94;
// bram[25447] = 78;
// bram[25448] = 62;
// bram[25449] = 48;
// bram[25450] = 35;
// bram[25451] = 24;
// bram[25452] = 15;
// bram[25453] = 7;
// bram[25454] = 2;
// bram[25455] = 0;
// bram[25456] = 0;
// bram[25457] = 2;
// bram[25458] = 6;
// bram[25459] = 13;
// bram[25460] = 22;
// bram[25461] = 33;
// bram[25462] = 45;
// bram[25463] = 60;
// bram[25464] = 75;
// bram[25465] = 91;
// bram[25466] = 108;
// bram[25467] = 126;
// bram[25468] = 143;
// bram[25469] = 160;
// bram[25470] = 176;
// bram[25471] = 192;
// bram[25472] = 206;
// bram[25473] = 219;
// bram[25474] = 230;
// bram[25475] = 239;
// bram[25476] = 246;
// bram[25477] = 251;
// bram[25478] = 253;
// bram[25479] = 253;
// bram[25480] = 251;
// bram[25481] = 246;
// bram[25482] = 239;
// bram[25483] = 230;
// bram[25484] = 219;
// bram[25485] = 206;
// bram[25486] = 192;
// bram[25487] = 177;
// bram[25488] = 160;
// bram[25489] = 143;
// bram[25490] = 126;
// bram[25491] = 109;
// bram[25492] = 92;
// bram[25493] = 75;
// bram[25494] = 60;
// bram[25495] = 46;
// bram[25496] = 33;
// bram[25497] = 22;
// bram[25498] = 13;
// bram[25499] = 6;
// bram[25500] = 2;
// bram[25501] = 0;
// bram[25502] = 0;
// bram[25503] = 2;
// bram[25504] = 7;
// bram[25505] = 14;
// bram[25506] = 24;
// bram[25507] = 35;
// bram[25508] = 48;
// bram[25509] = 62;
// bram[25510] = 77;
// bram[25511] = 94;
// bram[25512] = 111;
// bram[25513] = 128;
// bram[25514] = 146;
// bram[25515] = 163;
// bram[25516] = 179;
// bram[25517] = 194;
// bram[25518] = 208;
// bram[25519] = 221;
// bram[25520] = 232;
// bram[25521] = 240;
// bram[25522] = 247;
// bram[25523] = 251;
// bram[25524] = 253;
// bram[25525] = 253;
// bram[25526] = 250;
// bram[25527] = 245;
// bram[25528] = 238;
// bram[25529] = 229;
// bram[25530] = 217;
// bram[25531] = 204;
// bram[25532] = 190;
// bram[25533] = 174;
// bram[25534] = 158;
// bram[25535] = 141;
// bram[25536] = 123;
// bram[25537] = 106;
// bram[25538] = 89;
// bram[25539] = 73;
// bram[25540] = 58;
// bram[25541] = 44;
// bram[25542] = 31;
// bram[25543] = 21;
// bram[25544] = 12;
// bram[25545] = 6;
// bram[25546] = 1;
// bram[25547] = 0;
// bram[25548] = 0;
// bram[25549] = 3;
// bram[25550] = 8;
// bram[25551] = 16;
// bram[25552] = 25;
// bram[25553] = 37;
// bram[25554] = 50;
// bram[25555] = 64;
// bram[25556] = 80;
// bram[25557] = 97;
// bram[25558] = 114;
// bram[25559] = 131;
// bram[25560] = 148;
// bram[25561] = 165;
// bram[25562] = 181;
// bram[25563] = 197;
// bram[25564] = 210;
// bram[25565] = 223;
// bram[25566] = 233;
// bram[25567] = 241;
// bram[25568] = 248;
// bram[25569] = 252;
// bram[25570] = 253;
// bram[25571] = 253;
// bram[25572] = 250;
// bram[25573] = 244;
// bram[25574] = 237;
// bram[25575] = 227;
// bram[25576] = 215;
// bram[25577] = 202;
// bram[25578] = 188;
// bram[25579] = 172;
// bram[25580] = 155;
// bram[25581] = 138;
// bram[25582] = 121;
// bram[25583] = 103;
// bram[25584] = 86;
// bram[25585] = 70;
// bram[25586] = 55;
// bram[25587] = 42;
// bram[25588] = 30;
// bram[25589] = 19;
// bram[25590] = 11;
// bram[25591] = 5;
// bram[25592] = 1;
// bram[25593] = 0;
// bram[25594] = 0;
// bram[25595] = 4;
// bram[25596] = 9;
// bram[25597] = 17;
// bram[25598] = 27;
// bram[25599] = 39;
// bram[25600] = 52;
// bram[25601] = 67;
// bram[25602] = 82;
// bram[25603] = 99;
// bram[25604] = 116;
// bram[25605] = 134;
// bram[25606] = 151;
// bram[25607] = 168;
// bram[25608] = 184;
// bram[25609] = 199;
// bram[25610] = 212;
// bram[25611] = 224;
// bram[25612] = 234;
// bram[25613] = 243;
// bram[25614] = 249;
// bram[25615] = 252;
// bram[25616] = 253;
// bram[25617] = 252;
// bram[25618] = 249;
// bram[25619] = 243;
// bram[25620] = 235;
// bram[25621] = 225;
// bram[25622] = 214;
// bram[25623] = 200;
// bram[25624] = 185;
// bram[25625] = 169;
// bram[25626] = 153;
// bram[25627] = 135;
// bram[25628] = 118;
// bram[25629] = 101;
// bram[25630] = 84;
// bram[25631] = 68;
// bram[25632] = 53;
// bram[25633] = 40;
// bram[25634] = 28;
// bram[25635] = 18;
// bram[25636] = 10;
// bram[25637] = 4;
// bram[25638] = 1;
// bram[25639] = 0;
// bram[25640] = 1;
// bram[25641] = 4;
// bram[25642] = 10;
// bram[25643] = 18;
// bram[25644] = 29;
// bram[25645] = 40;
// bram[25646] = 54;
// bram[25647] = 69;
// bram[25648] = 85;
// bram[25649] = 102;
// bram[25650] = 119;
// bram[25651] = 136;
// bram[25652] = 154;
// bram[25653] = 170;
// bram[25654] = 186;
// bram[25655] = 201;
// bram[25656] = 214;
// bram[25657] = 226;
// bram[25658] = 236;
// bram[25659] = 244;
// bram[25660] = 249;
// bram[25661] = 253;
// bram[25662] = 253;
// bram[25663] = 252;
// bram[25664] = 248;
// bram[25665] = 242;
// bram[25666] = 234;
// bram[25667] = 224;
// bram[25668] = 212;
// bram[25669] = 198;
// bram[25670] = 183;
// bram[25671] = 167;
// bram[25672] = 150;
// bram[25673] = 133;
// bram[25674] = 115;
// bram[25675] = 98;
// bram[25676] = 81;
// bram[25677] = 66;
// bram[25678] = 51;
// bram[25679] = 38;
// bram[25680] = 26;
// bram[25681] = 16;
// bram[25682] = 9;
// bram[25683] = 3;
// bram[25684] = 0;
// bram[25685] = 0;
// bram[25686] = 1;
// bram[25687] = 5;
// bram[25688] = 11;
// bram[25689] = 20;
// bram[25690] = 30;
// bram[25691] = 42;
// bram[25692] = 56;
// bram[25693] = 71;
// bram[25694] = 88;
// bram[25695] = 104;
// bram[25696] = 122;
// bram[25697] = 139;
// bram[25698] = 156;
// bram[25699] = 173;
// bram[25700] = 189;
// bram[25701] = 203;
// bram[25702] = 216;
// bram[25703] = 228;
// bram[25704] = 237;
// bram[25705] = 245;
// bram[25706] = 250;
// bram[25707] = 253;
// bram[25708] = 253;
// bram[25709] = 252;
// bram[25710] = 247;
// bram[25711] = 241;
// bram[25712] = 232;
// bram[25713] = 222;
// bram[25714] = 210;
// bram[25715] = 196;
// bram[25716] = 180;
// bram[25717] = 164;
// bram[25718] = 147;
// bram[25719] = 130;
// bram[25720] = 113;
// bram[25721] = 95;
// bram[25722] = 79;
// bram[25723] = 63;
// bram[25724] = 49;
// bram[25725] = 36;
// bram[25726] = 25;
// bram[25727] = 15;
// bram[25728] = 8;
// bram[25729] = 3;
// bram[25730] = 0;
// bram[25731] = 0;
// bram[25732] = 2;
// bram[25733] = 6;
// bram[25734] = 13;
// bram[25735] = 21;
// bram[25736] = 32;
// bram[25737] = 45;
// bram[25738] = 59;
// bram[25739] = 74;
// bram[25740] = 90;
// bram[25741] = 107;
// bram[25742] = 124;
// bram[25743] = 142;
// bram[25744] = 159;
// bram[25745] = 175;
// bram[25746] = 191;
// bram[25747] = 205;
// bram[25748] = 218;
// bram[25749] = 229;
// bram[25750] = 239;
// bram[25751] = 246;
// bram[25752] = 251;
// bram[25753] = 253;
// bram[25754] = 253;
// bram[25755] = 251;
// bram[25756] = 247;
// bram[25757] = 240;
// bram[25758] = 231;
// bram[25759] = 220;
// bram[25760] = 207;
// bram[25761] = 193;
// bram[25762] = 178;
// bram[25763] = 162;
// bram[25764] = 145;
// bram[25765] = 127;
// bram[25766] = 110;
// bram[25767] = 93;
// bram[25768] = 76;
// bram[25769] = 61;
// bram[25770] = 47;
// bram[25771] = 34;
// bram[25772] = 23;
// bram[25773] = 14;
// bram[25774] = 7;
// bram[25775] = 2;
// bram[25776] = 0;
// bram[25777] = 0;
// bram[25778] = 2;
// bram[25779] = 7;
// bram[25780] = 14;
// bram[25781] = 23;
// bram[25782] = 34;
// bram[25783] = 47;
// bram[25784] = 61;
// bram[25785] = 76;
// bram[25786] = 93;
// bram[25787] = 110;
// bram[25788] = 127;
// bram[25789] = 144;
// bram[25790] = 161;
// bram[25791] = 178;
// bram[25792] = 193;
// bram[25793] = 207;
// bram[25794] = 220;
// bram[25795] = 231;
// bram[25796] = 240;
// bram[25797] = 247;
// bram[25798] = 251;
// bram[25799] = 253;
// bram[25800] = 253;
// bram[25801] = 251;
// bram[25802] = 246;
// bram[25803] = 239;
// bram[25804] = 229;
// bram[25805] = 218;
// bram[25806] = 205;
// bram[25807] = 191;
// bram[25808] = 175;
// bram[25809] = 159;
// bram[25810] = 142;
// bram[25811] = 125;
// bram[25812] = 107;
// bram[25813] = 90;
// bram[25814] = 74;
// bram[25815] = 59;
// bram[25816] = 45;
// bram[25817] = 32;
// bram[25818] = 21;
// bram[25819] = 13;
// bram[25820] = 6;
// bram[25821] = 2;
// bram[25822] = 0;
// bram[25823] = 0;
// bram[25824] = 3;
// bram[25825] = 8;
// bram[25826] = 15;
// bram[25827] = 24;
// bram[25828] = 36;
// bram[25829] = 49;
// bram[25830] = 63;
// bram[25831] = 79;
// bram[25832] = 95;
// bram[25833] = 112;
// bram[25834] = 130;
// bram[25835] = 147;
// bram[25836] = 164;
// bram[25837] = 180;
// bram[25838] = 195;
// bram[25839] = 209;
// bram[25840] = 222;
// bram[25841] = 232;
// bram[25842] = 241;
// bram[25843] = 247;
// bram[25844] = 252;
// bram[25845] = 253;
// bram[25846] = 253;
// bram[25847] = 250;
// bram[25848] = 245;
// bram[25849] = 237;
// bram[25850] = 228;
// bram[25851] = 216;
// bram[25852] = 203;
// bram[25853] = 189;
// bram[25854] = 173;
// bram[25855] = 156;
// bram[25856] = 139;
// bram[25857] = 122;
// bram[25858] = 105;
// bram[25859] = 88;
// bram[25860] = 72;
// bram[25861] = 56;
// bram[25862] = 43;
// bram[25863] = 30;
// bram[25864] = 20;
// bram[25865] = 11;
// bram[25866] = 5;
// bram[25867] = 1;
// bram[25868] = 0;
// bram[25869] = 0;
// bram[25870] = 3;
// bram[25871] = 9;
// bram[25872] = 16;
// bram[25873] = 26;
// bram[25874] = 38;
// bram[25875] = 51;
// bram[25876] = 65;
// bram[25877] = 81;
// bram[25878] = 98;
// bram[25879] = 115;
// bram[25880] = 132;
// bram[25881] = 150;
// bram[25882] = 167;
// bram[25883] = 183;
// bram[25884] = 198;
// bram[25885] = 211;
// bram[25886] = 224;
// bram[25887] = 234;
// bram[25888] = 242;
// bram[25889] = 248;
// bram[25890] = 252;
// bram[25891] = 253;
// bram[25892] = 253;
// bram[25893] = 249;
// bram[25894] = 244;
// bram[25895] = 236;
// bram[25896] = 226;
// bram[25897] = 214;
// bram[25898] = 201;
// bram[25899] = 186;
// bram[25900] = 170;
// bram[25901] = 154;
// bram[25902] = 137;
// bram[25903] = 119;
// bram[25904] = 102;
// bram[25905] = 85;
// bram[25906] = 69;
// bram[25907] = 54;
// bram[25908] = 41;
// bram[25909] = 29;
// bram[25910] = 18;
// bram[25911] = 10;
// bram[25912] = 4;
// bram[25913] = 1;
// bram[25914] = 0;
// bram[25915] = 1;
// bram[25916] = 4;
// bram[25917] = 10;
// bram[25918] = 18;
// bram[25919] = 28;
// bram[25920] = 40;
// bram[25921] = 53;
// bram[25922] = 68;
// bram[25923] = 84;
// bram[25924] = 101;
// bram[25925] = 118;
// bram[25926] = 135;
// bram[25927] = 152;
// bram[25928] = 169;
// bram[25929] = 185;
// bram[25930] = 200;
// bram[25931] = 213;
// bram[25932] = 225;
// bram[25933] = 235;
// bram[25934] = 243;
// bram[25935] = 249;
// bram[25936] = 252;
// bram[25937] = 253;
// bram[25938] = 252;
// bram[25939] = 249;
// bram[25940] = 243;
// bram[25941] = 235;
// bram[25942] = 224;
// bram[25943] = 212;
// bram[25944] = 199;
// bram[25945] = 184;
// bram[25946] = 168;
// bram[25947] = 151;
// bram[25948] = 134;
// bram[25949] = 116;
// bram[25950] = 99;
// bram[25951] = 83;
// bram[25952] = 67;
// bram[25953] = 52;
// bram[25954] = 39;
// bram[25955] = 27;
// bram[25956] = 17;
// bram[25957] = 9;
// bram[25958] = 4;
// bram[25959] = 0;
// bram[25960] = 0;
// bram[25961] = 1;
// bram[25962] = 5;
// bram[25963] = 11;
// bram[25964] = 19;
// bram[25965] = 29;
// bram[25966] = 42;
// bram[25967] = 55;
// bram[25968] = 70;
// bram[25969] = 86;
// bram[25970] = 103;
// bram[25971] = 120;
// bram[25972] = 138;
// bram[25973] = 155;
// bram[25974] = 172;
// bram[25975] = 187;
// bram[25976] = 202;
// bram[25977] = 215;
// bram[25978] = 227;
// bram[25979] = 237;
// bram[25980] = 244;
// bram[25981] = 250;
// bram[25982] = 253;
// bram[25983] = 253;
// bram[25984] = 252;
// bram[25985] = 248;
// bram[25986] = 242;
// bram[25987] = 233;
// bram[25988] = 223;
// bram[25989] = 210;
// bram[25990] = 197;
// bram[25991] = 182;
// bram[25992] = 165;
// bram[25993] = 148;
// bram[25994] = 131;
// bram[25995] = 114;
// bram[25996] = 97;
// bram[25997] = 80;
// bram[25998] = 64;
// bram[25999] = 50;
// bram[26000] = 37;
// bram[26001] = 25;
// bram[26002] = 16;
// bram[26003] = 8;
// bram[26004] = 3;
// bram[26005] = 0;
// bram[26006] = 0;
// bram[26007] = 1;
// bram[26008] = 6;
// bram[26009] = 12;
// bram[26010] = 21;
// bram[26011] = 31;
// bram[26012] = 44;
// bram[26013] = 57;
// bram[26014] = 73;
// bram[26015] = 89;
// bram[26016] = 106;
// bram[26017] = 123;
// bram[26018] = 141;
// bram[26019] = 158;
// bram[26020] = 174;
// bram[26021] = 190;
// bram[26022] = 204;
// bram[26023] = 217;
// bram[26024] = 229;
// bram[26025] = 238;
// bram[26026] = 245;
// bram[26027] = 250;
// bram[26028] = 253;
// bram[26029] = 253;
// bram[26030] = 251;
// bram[26031] = 247;
// bram[26032] = 240;
// bram[26033] = 232;
// bram[26034] = 221;
// bram[26035] = 208;
// bram[26036] = 194;
// bram[26037] = 179;
// bram[26038] = 163;
// bram[26039] = 146;
// bram[26040] = 128;
// bram[26041] = 111;
// bram[26042] = 94;
// bram[26043] = 78;
// bram[26044] = 62;
// bram[26045] = 48;
// bram[26046] = 35;
// bram[26047] = 24;
// bram[26048] = 14;
// bram[26049] = 7;
// bram[26050] = 2;
// bram[26051] = 0;
// bram[26052] = 0;
// bram[26053] = 2;
// bram[26054] = 6;
// bram[26055] = 13;
// bram[26056] = 22;
// bram[26057] = 33;
// bram[26058] = 46;
// bram[26059] = 60;
// bram[26060] = 75;
// bram[26061] = 91;
// bram[26062] = 109;
// bram[26063] = 126;
// bram[26064] = 143;
// bram[26065] = 160;
// bram[26066] = 177;
// bram[26067] = 192;
// bram[26068] = 206;
// bram[26069] = 219;
// bram[26070] = 230;
// bram[26071] = 239;
// bram[26072] = 246;
// bram[26073] = 251;
// bram[26074] = 253;
// bram[26075] = 253;
// bram[26076] = 251;
// bram[26077] = 246;
// bram[26078] = 239;
// bram[26079] = 230;
// bram[26080] = 219;
// bram[26081] = 206;
// bram[26082] = 192;
// bram[26083] = 177;
// bram[26084] = 160;
// bram[26085] = 143;
// bram[26086] = 126;
// bram[26087] = 108;
// bram[26088] = 91;
// bram[26089] = 75;
// bram[26090] = 60;
// bram[26091] = 46;
// bram[26092] = 33;
// bram[26093] = 22;
// bram[26094] = 13;
// bram[26095] = 6;
// bram[26096] = 2;
// bram[26097] = 0;
// bram[26098] = 0;
// bram[26099] = 2;
// bram[26100] = 7;
// bram[26101] = 14;
// bram[26102] = 24;
// bram[26103] = 35;
// bram[26104] = 48;
// bram[26105] = 62;
// bram[26106] = 78;
// bram[26107] = 94;
// bram[26108] = 111;
// bram[26109] = 129;
// bram[26110] = 146;
// bram[26111] = 163;
// bram[26112] = 179;
// bram[26113] = 194;
// bram[26114] = 208;
// bram[26115] = 221;
// bram[26116] = 232;
// bram[26117] = 240;
// bram[26118] = 247;
// bram[26119] = 251;
// bram[26120] = 253;
// bram[26121] = 253;
// bram[26122] = 250;
// bram[26123] = 245;
// bram[26124] = 238;
// bram[26125] = 229;
// bram[26126] = 217;
// bram[26127] = 204;
// bram[26128] = 190;
// bram[26129] = 174;
// bram[26130] = 158;
// bram[26131] = 140;
// bram[26132] = 123;
// bram[26133] = 106;
// bram[26134] = 89;
// bram[26135] = 73;
// bram[26136] = 57;
// bram[26137] = 44;
// bram[26138] = 31;
// bram[26139] = 21;
// bram[26140] = 12;
// bram[26141] = 6;
// bram[26142] = 1;
// bram[26143] = 0;
// bram[26144] = 0;
// bram[26145] = 3;
// bram[26146] = 8;
// bram[26147] = 16;
// bram[26148] = 25;
// bram[26149] = 37;
// bram[26150] = 50;
// bram[26151] = 64;
// bram[26152] = 80;
// bram[26153] = 97;
// bram[26154] = 114;
// bram[26155] = 131;
// bram[26156] = 149;
// bram[26157] = 165;
// bram[26158] = 182;
// bram[26159] = 197;
// bram[26160] = 210;
// bram[26161] = 223;
// bram[26162] = 233;
// bram[26163] = 242;
// bram[26164] = 248;
// bram[26165] = 252;
// bram[26166] = 253;
// bram[26167] = 253;
// bram[26168] = 250;
// bram[26169] = 244;
// bram[26170] = 237;
// bram[26171] = 227;
// bram[26172] = 215;
// bram[26173] = 202;
// bram[26174] = 187;
// bram[26175] = 172;
// bram[26176] = 155;
// bram[26177] = 138;
// bram[26178] = 120;
// bram[26179] = 103;
// bram[26180] = 86;
// bram[26181] = 70;
// bram[26182] = 55;
// bram[26183] = 42;
// bram[26184] = 29;
// bram[26185] = 19;
// bram[26186] = 11;
// bram[26187] = 5;
// bram[26188] = 1;
// bram[26189] = 0;
// bram[26190] = 0;
// bram[26191] = 4;
// bram[26192] = 9;
// bram[26193] = 17;
// bram[26194] = 27;
// bram[26195] = 39;
// bram[26196] = 52;
// bram[26197] = 67;
// bram[26198] = 83;
// bram[26199] = 99;
// bram[26200] = 117;
// bram[26201] = 134;
// bram[26202] = 151;
// bram[26203] = 168;
// bram[26204] = 184;
// bram[26205] = 199;
// bram[26206] = 212;
// bram[26207] = 224;
// bram[26208] = 235;
// bram[26209] = 243;
// bram[26210] = 249;
// bram[26211] = 252;
// bram[26212] = 253;
// bram[26213] = 252;
// bram[26214] = 249;
// bram[26215] = 243;
// bram[26216] = 235;
// bram[26217] = 225;
// bram[26218] = 213;
// bram[26219] = 200;
// bram[26220] = 185;
// bram[26221] = 169;
// bram[26222] = 152;
// bram[26223] = 135;
// bram[26224] = 118;
// bram[26225] = 101;
// bram[26226] = 84;
// bram[26227] = 68;
// bram[26228] = 53;
// bram[26229] = 40;
// bram[26230] = 28;
// bram[26231] = 18;
// bram[26232] = 10;
// bram[26233] = 4;
// bram[26234] = 1;
// bram[26235] = 0;
// bram[26236] = 1;
// bram[26237] = 4;
// bram[26238] = 10;
// bram[26239] = 19;
// bram[26240] = 29;
// bram[26241] = 41;
// bram[26242] = 54;
// bram[26243] = 69;
// bram[26244] = 85;
// bram[26245] = 102;
// bram[26246] = 119;
// bram[26247] = 137;
// bram[26248] = 154;
// bram[26249] = 171;
// bram[26250] = 186;
// bram[26251] = 201;
// bram[26252] = 214;
// bram[26253] = 226;
// bram[26254] = 236;
// bram[26255] = 244;
// bram[26256] = 249;
// bram[26257] = 253;
// bram[26258] = 253;
// bram[26259] = 252;
// bram[26260] = 248;
// bram[26261] = 242;
// bram[26262] = 234;
// bram[26263] = 223;
// bram[26264] = 211;
// bram[26265] = 198;
// bram[26266] = 183;
// bram[26267] = 167;
// bram[26268] = 150;
// bram[26269] = 132;
// bram[26270] = 115;
// bram[26271] = 98;
// bram[26272] = 81;
// bram[26273] = 65;
// bram[26274] = 51;
// bram[26275] = 38;
// bram[26276] = 26;
// bram[26277] = 16;
// bram[26278] = 9;
// bram[26279] = 3;
// bram[26280] = 0;
// bram[26281] = 0;
// bram[26282] = 1;
// bram[26283] = 5;
// bram[26284] = 12;
// bram[26285] = 20;
// bram[26286] = 30;
// bram[26287] = 43;
// bram[26288] = 56;
// bram[26289] = 72;
// bram[26290] = 88;
// bram[26291] = 105;
// bram[26292] = 122;
// bram[26293] = 139;
// bram[26294] = 156;
// bram[26295] = 173;
// bram[26296] = 189;
// bram[26297] = 203;
// bram[26298] = 216;
// bram[26299] = 228;
// bram[26300] = 237;
// bram[26301] = 245;
// bram[26302] = 250;
// bram[26303] = 253;
// bram[26304] = 253;
// bram[26305] = 252;
// bram[26306] = 247;
// bram[26307] = 241;
// bram[26308] = 232;
// bram[26309] = 222;
// bram[26310] = 209;
// bram[26311] = 195;
// bram[26312] = 180;
// bram[26313] = 164;
// bram[26314] = 147;
// bram[26315] = 130;
// bram[26316] = 112;
// bram[26317] = 95;
// bram[26318] = 79;
// bram[26319] = 63;
// bram[26320] = 49;
// bram[26321] = 36;
// bram[26322] = 24;
// bram[26323] = 15;
// bram[26324] = 8;
// bram[26325] = 3;
// bram[26326] = 0;
// bram[26327] = 0;
// bram[26328] = 2;
// bram[26329] = 6;
// bram[26330] = 13;
// bram[26331] = 21;
// bram[26332] = 32;
// bram[26333] = 45;
// bram[26334] = 59;
// bram[26335] = 74;
// bram[26336] = 90;
// bram[26337] = 107;
// bram[26338] = 125;
// bram[26339] = 142;
// bram[26340] = 159;
// bram[26341] = 176;
// bram[26342] = 191;
// bram[26343] = 205;
// bram[26344] = 218;
// bram[26345] = 229;
// bram[26346] = 239;
// bram[26347] = 246;
// bram[26348] = 251;
// bram[26349] = 253;
// bram[26350] = 253;
// bram[26351] = 251;
// bram[26352] = 247;
// bram[26353] = 240;
// bram[26354] = 231;
// bram[26355] = 220;
// bram[26356] = 207;
// bram[26357] = 193;
// bram[26358] = 178;
// bram[26359] = 161;
// bram[26360] = 144;
// bram[26361] = 127;
// bram[26362] = 110;
// bram[26363] = 93;
// bram[26364] = 76;
// bram[26365] = 61;
// bram[26366] = 47;
// bram[26367] = 34;
// bram[26368] = 23;
// bram[26369] = 14;
// bram[26370] = 7;
// bram[26371] = 2;
// bram[26372] = 0;
// bram[26373] = 0;
// bram[26374] = 2;
// bram[26375] = 7;
// bram[26376] = 14;
// bram[26377] = 23;
// bram[26378] = 34;
// bram[26379] = 47;
// bram[26380] = 61;
// bram[26381] = 76;
// bram[26382] = 93;
// bram[26383] = 110;
// bram[26384] = 127;
// bram[26385] = 145;
// bram[26386] = 162;
// bram[26387] = 178;
// bram[26388] = 193;
// bram[26389] = 207;
// bram[26390] = 220;
// bram[26391] = 231;
// bram[26392] = 240;
// bram[26393] = 247;
// bram[26394] = 251;
// bram[26395] = 253;
// bram[26396] = 253;
// bram[26397] = 251;
// bram[26398] = 246;
// bram[26399] = 238;
// bram[26400] = 229;
// bram[26401] = 218;
// bram[26402] = 205;
// bram[26403] = 191;
// bram[26404] = 175;
// bram[26405] = 159;
// bram[26406] = 142;
// bram[26407] = 124;
// bram[26408] = 107;
// bram[26409] = 90;
// bram[26410] = 74;
// bram[26411] = 58;
// bram[26412] = 44;
// bram[26413] = 32;
// bram[26414] = 21;
// bram[26415] = 13;
// bram[26416] = 6;
// bram[26417] = 2;
// bram[26418] = 0;
// bram[26419] = 0;
// bram[26420] = 3;
// bram[26421] = 8;
// bram[26422] = 15;
// bram[26423] = 25;
// bram[26424] = 36;
// bram[26425] = 49;
// bram[26426] = 63;
// bram[26427] = 79;
// bram[26428] = 95;
// bram[26429] = 113;
// bram[26430] = 130;
// bram[26431] = 147;
// bram[26432] = 164;
// bram[26433] = 180;
// bram[26434] = 196;
// bram[26435] = 210;
// bram[26436] = 222;
// bram[26437] = 232;
// bram[26438] = 241;
// bram[26439] = 247;
// bram[26440] = 252;
// bram[26441] = 253;
// bram[26442] = 253;
// bram[26443] = 250;
// bram[26444] = 245;
// bram[26445] = 237;
// bram[26446] = 228;
// bram[26447] = 216;
// bram[26448] = 203;
// bram[26449] = 189;
// bram[26450] = 173;
// bram[26451] = 156;
// bram[26452] = 139;
// bram[26453] = 122;
// bram[26454] = 104;
// bram[26455] = 87;
// bram[26456] = 71;
// bram[26457] = 56;
// bram[26458] = 42;
// bram[26459] = 30;
// bram[26460] = 20;
// bram[26461] = 11;
// bram[26462] = 5;
// bram[26463] = 1;
// bram[26464] = 0;
// bram[26465] = 0;
// bram[26466] = 3;
// bram[26467] = 9;
// bram[26468] = 16;
// bram[26469] = 26;
// bram[26470] = 38;
// bram[26471] = 51;
// bram[26472] = 66;
// bram[26473] = 81;
// bram[26474] = 98;
// bram[26475] = 115;
// bram[26476] = 133;
// bram[26477] = 150;
// bram[26478] = 167;
// bram[26479] = 183;
// bram[26480] = 198;
// bram[26481] = 212;
// bram[26482] = 224;
// bram[26483] = 234;
// bram[26484] = 242;
// bram[26485] = 248;
// bram[26486] = 252;
// bram[26487] = 253;
// bram[26488] = 253;
// bram[26489] = 249;
// bram[26490] = 244;
// bram[26491] = 236;
// bram[26492] = 226;
// bram[26493] = 214;
// bram[26494] = 201;
// bram[26495] = 186;
// bram[26496] = 170;
// bram[26497] = 154;
// bram[26498] = 136;
// bram[26499] = 119;
// bram[26500] = 102;
// bram[26501] = 85;
// bram[26502] = 69;
// bram[26503] = 54;
// bram[26504] = 40;
// bram[26505] = 28;
// bram[26506] = 18;
// bram[26507] = 10;
// bram[26508] = 4;
// bram[26509] = 1;
// bram[26510] = 0;
// bram[26511] = 1;
// bram[26512] = 4;
// bram[26513] = 10;
// bram[26514] = 18;
// bram[26515] = 28;
// bram[26516] = 40;
// bram[26517] = 53;
// bram[26518] = 68;
// bram[26519] = 84;
// bram[26520] = 101;
// bram[26521] = 118;
// bram[26522] = 135;
// bram[26523] = 153;
// bram[26524] = 169;
// bram[26525] = 185;
// bram[26526] = 200;
// bram[26527] = 214;
// bram[26528] = 225;
// bram[26529] = 235;
// bram[26530] = 243;
// bram[26531] = 249;
// bram[26532] = 252;
// bram[26533] = 253;
// bram[26534] = 252;
// bram[26535] = 249;
// bram[26536] = 243;
// bram[26537] = 234;
// bram[26538] = 224;
// bram[26539] = 212;
// bram[26540] = 199;
// bram[26541] = 184;
// bram[26542] = 168;
// bram[26543] = 151;
// bram[26544] = 134;
// bram[26545] = 116;
// bram[26546] = 99;
// bram[26547] = 82;
// bram[26548] = 67;
// bram[26549] = 52;
// bram[26550] = 38;
// bram[26551] = 27;
// bram[26552] = 17;
// bram[26553] = 9;
// bram[26554] = 4;
// bram[26555] = 0;
// bram[26556] = 0;
// bram[26557] = 1;
// bram[26558] = 5;
// bram[26559] = 11;
// bram[26560] = 19;
// bram[26561] = 30;
// bram[26562] = 42;
// bram[26563] = 55;
// bram[26564] = 70;
// bram[26565] = 87;
// bram[26566] = 103;
// bram[26567] = 121;
// bram[26568] = 138;
// bram[26569] = 155;
// bram[26570] = 172;
// bram[26571] = 188;
// bram[26572] = 202;
// bram[26573] = 215;
// bram[26574] = 227;
// bram[26575] = 237;
// bram[26576] = 244;
// bram[26577] = 250;
// bram[26578] = 253;
// bram[26579] = 253;
// bram[26580] = 252;
// bram[26581] = 248;
// bram[26582] = 241;
// bram[26583] = 233;
// bram[26584] = 223;
// bram[26585] = 210;
// bram[26586] = 196;
// bram[26587] = 181;
// bram[26588] = 165;
// bram[26589] = 148;
// bram[26590] = 131;
// bram[26591] = 114;
// bram[26592] = 96;
// bram[26593] = 80;
// bram[26594] = 64;
// bram[26595] = 50;
// bram[26596] = 37;
// bram[26597] = 25;
// bram[26598] = 16;
// bram[26599] = 8;
// bram[26600] = 3;
// bram[26601] = 0;
// bram[26602] = 0;
// bram[26603] = 1;
// bram[26604] = 6;
// bram[26605] = 12;
// bram[26606] = 21;
// bram[26607] = 31;
// bram[26608] = 44;
// bram[26609] = 58;
// bram[26610] = 73;
// bram[26611] = 89;
// bram[26612] = 106;
// bram[26613] = 123;
// bram[26614] = 141;
// bram[26615] = 158;
// bram[26616] = 174;
// bram[26617] = 190;
// bram[26618] = 204;
// bram[26619] = 217;
// bram[26620] = 229;
// bram[26621] = 238;
// bram[26622] = 245;
// bram[26623] = 250;
// bram[26624] = 253;
// bram[26625] = 253;
// bram[26626] = 251;
// bram[26627] = 247;
// bram[26628] = 240;
// bram[26629] = 232;
// bram[26630] = 221;
// bram[26631] = 208;
// bram[26632] = 194;
// bram[26633] = 179;
// bram[26634] = 163;
// bram[26635] = 146;
// bram[26636] = 128;
// bram[26637] = 111;
// bram[26638] = 94;
// bram[26639] = 77;
// bram[26640] = 62;
// bram[26641] = 48;
// bram[26642] = 35;
// bram[26643] = 24;
// bram[26644] = 14;
// bram[26645] = 7;
// bram[26646] = 2;
// bram[26647] = 0;
// bram[26648] = 0;
// bram[26649] = 2;
// bram[26650] = 7;
// bram[26651] = 13;
// bram[26652] = 22;
// bram[26653] = 33;
// bram[26654] = 46;
// bram[26655] = 60;
// bram[26656] = 75;
// bram[26657] = 92;
// bram[26658] = 109;
// bram[26659] = 126;
// bram[26660] = 143;
// bram[26661] = 160;
// bram[26662] = 177;
// bram[26663] = 192;
// bram[26664] = 207;
// bram[26665] = 219;
// bram[26666] = 230;
// bram[26667] = 239;
// bram[26668] = 246;
// bram[26669] = 251;
// bram[26670] = 253;
// bram[26671] = 253;
// bram[26672] = 251;
// bram[26673] = 246;
// bram[26674] = 239;
// bram[26675] = 230;
// bram[26676] = 219;
// bram[26677] = 206;
// bram[26678] = 192;
// bram[26679] = 176;
// bram[26680] = 160;
// bram[26681] = 143;
// bram[26682] = 126;
// bram[26683] = 108;
// bram[26684] = 91;
// bram[26685] = 75;
// bram[26686] = 60;
// bram[26687] = 45;
// bram[26688] = 33;
// bram[26689] = 22;
// bram[26690] = 13;
// bram[26691] = 6;
// bram[26692] = 2;
// bram[26693] = 0;
// bram[26694] = 0;
// bram[26695] = 3;
// bram[26696] = 7;
// bram[26697] = 15;
// bram[26698] = 24;
// bram[26699] = 35;
// bram[26700] = 48;
// bram[26701] = 62;
// bram[26702] = 78;
// bram[26703] = 94;
// bram[26704] = 111;
// bram[26705] = 129;
// bram[26706] = 146;
// bram[26707] = 163;
// bram[26708] = 179;
// bram[26709] = 195;
// bram[26710] = 209;
// bram[26711] = 221;
// bram[26712] = 232;
// bram[26713] = 240;
// bram[26714] = 247;
// bram[26715] = 251;
// bram[26716] = 253;
// bram[26717] = 253;
// bram[26718] = 250;
// bram[26719] = 245;
// bram[26720] = 238;
// bram[26721] = 228;
// bram[26722] = 217;
// bram[26723] = 204;
// bram[26724] = 190;
// bram[26725] = 174;
// bram[26726] = 157;
// bram[26727] = 140;
// bram[26728] = 123;
// bram[26729] = 106;
// bram[26730] = 89;
// bram[26731] = 72;
// bram[26732] = 57;
// bram[26733] = 43;
// bram[26734] = 31;
// bram[26735] = 20;
// bram[26736] = 12;
// bram[26737] = 6;
// bram[26738] = 1;
// bram[26739] = 0;
// bram[26740] = 0;
// bram[26741] = 3;
// bram[26742] = 8;
// bram[26743] = 16;
// bram[26744] = 25;
// bram[26745] = 37;
// bram[26746] = 50;
// bram[26747] = 65;
// bram[26748] = 80;
// bram[26749] = 97;
// bram[26750] = 114;
// bram[26751] = 131;
// bram[26752] = 149;
// bram[26753] = 166;
// bram[26754] = 182;
// bram[26755] = 197;
// bram[26756] = 211;
// bram[26757] = 223;
// bram[26758] = 233;
// bram[26759] = 242;
// bram[26760] = 248;
// bram[26761] = 252;
// bram[26762] = 253;
// bram[26763] = 253;
// bram[26764] = 250;
// bram[26765] = 244;
// bram[26766] = 236;
// bram[26767] = 227;
// bram[26768] = 215;
// bram[26769] = 202;
// bram[26770] = 187;
// bram[26771] = 171;
// bram[26772] = 155;
// bram[26773] = 138;
// bram[26774] = 120;
// bram[26775] = 103;
// bram[26776] = 86;
// bram[26777] = 70;
// bram[26778] = 55;
// bram[26779] = 41;
// bram[26780] = 29;
// bram[26781] = 19;
// bram[26782] = 11;
// bram[26783] = 5;
// bram[26784] = 1;
// bram[26785] = 0;
// bram[26786] = 0;
// bram[26787] = 4;
// bram[26788] = 9;
// bram[26789] = 17;
// bram[26790] = 27;
// bram[26791] = 39;
// bram[26792] = 52;
// bram[26793] = 67;
// bram[26794] = 83;
// bram[26795] = 100;
// bram[26796] = 117;
// bram[26797] = 134;
// bram[26798] = 151;
// bram[26799] = 168;
// bram[26800] = 184;
// bram[26801] = 199;
// bram[26802] = 213;
// bram[26803] = 225;
// bram[26804] = 235;
// bram[26805] = 243;
// bram[26806] = 249;
// bram[26807] = 252;
// bram[26808] = 253;
// bram[26809] = 252;
// bram[26810] = 249;
// bram[26811] = 243;
// bram[26812] = 235;
// bram[26813] = 225;
// bram[26814] = 213;
// bram[26815] = 200;
// bram[26816] = 185;
// bram[26817] = 169;
// bram[26818] = 152;
// bram[26819] = 135;
// bram[26820] = 118;
// bram[26821] = 100;
// bram[26822] = 84;
// bram[26823] = 68;
// bram[26824] = 53;
// bram[26825] = 39;
// bram[26826] = 28;
// bram[26827] = 18;
// bram[26828] = 10;
// bram[26829] = 4;
// bram[26830] = 1;
// bram[26831] = 0;
// bram[26832] = 1;
// bram[26833] = 5;
// bram[26834] = 10;
// bram[26835] = 19;
// bram[26836] = 29;
// bram[26837] = 41;
// bram[26838] = 54;
// bram[26839] = 69;
// bram[26840] = 85;
// bram[26841] = 102;
// bram[26842] = 119;
// bram[26843] = 137;
// bram[26844] = 154;
// bram[26845] = 171;
// bram[26846] = 187;
// bram[26847] = 201;
// bram[26848] = 215;
// bram[26849] = 226;
// bram[26850] = 236;
// bram[26851] = 244;
// bram[26852] = 249;
// bram[26853] = 253;
// bram[26854] = 253;
// bram[26855] = 252;
// bram[26856] = 248;
// bram[26857] = 242;
// bram[26858] = 234;
// bram[26859] = 223;
// bram[26860] = 211;
// bram[26861] = 198;
// bram[26862] = 182;
// bram[26863] = 166;
// bram[26864] = 150;
// bram[26865] = 132;
// bram[26866] = 115;
// bram[26867] = 98;
// bram[26868] = 81;
// bram[26869] = 65;
// bram[26870] = 51;
// bram[26871] = 37;
// bram[26872] = 26;
// bram[26873] = 16;
// bram[26874] = 9;
// bram[26875] = 3;
// bram[26876] = 0;
// bram[26877] = 0;
// bram[26878] = 1;
// bram[26879] = 5;
// bram[26880] = 12;
// bram[26881] = 20;
// bram[26882] = 31;
// bram[26883] = 43;
// bram[26884] = 57;
// bram[26885] = 72;
// bram[26886] = 88;
// bram[26887] = 105;
// bram[26888] = 122;
// bram[26889] = 139;
// bram[26890] = 157;
// bram[26891] = 173;
// bram[26892] = 189;
// bram[26893] = 203;
// bram[26894] = 217;
// bram[26895] = 228;
// bram[26896] = 237;
// bram[26897] = 245;
// bram[26898] = 250;
// bram[26899] = 253;
// bram[26900] = 253;
// bram[26901] = 252;
// bram[26902] = 247;
// bram[26903] = 241;
// bram[26904] = 232;
// bram[26905] = 222;
// bram[26906] = 209;
// bram[26907] = 195;
// bram[26908] = 180;
// bram[26909] = 164;
// bram[26910] = 147;
// bram[26911] = 130;
// bram[26912] = 112;
// bram[26913] = 95;
// bram[26914] = 79;
// bram[26915] = 63;
// bram[26916] = 49;
// bram[26917] = 36;
// bram[26918] = 24;
// bram[26919] = 15;
// bram[26920] = 8;
// bram[26921] = 3;
// bram[26922] = 0;
// bram[26923] = 0;
// bram[26924] = 2;
// bram[26925] = 6;
// bram[26926] = 13;
// bram[26927] = 22;
// bram[26928] = 32;
// bram[26929] = 45;
// bram[26930] = 59;
// bram[26931] = 74;
// bram[26932] = 90;
// bram[26933] = 107;
// bram[26934] = 125;
// bram[26935] = 142;
// bram[26936] = 159;
// bram[26937] = 176;
// bram[26938] = 191;
// bram[26939] = 206;
// bram[26940] = 218;
// bram[26941] = 230;
// bram[26942] = 239;
// bram[26943] = 246;
// bram[26944] = 251;
// bram[26945] = 253;
// bram[26946] = 253;
// bram[26947] = 251;
// bram[26948] = 246;
// bram[26949] = 240;
// bram[26950] = 231;
// bram[26951] = 220;
// bram[26952] = 207;
// bram[26953] = 193;
// bram[26954] = 178;
// bram[26955] = 161;
// bram[26956] = 144;
// bram[26957] = 127;
// bram[26958] = 109;
// bram[26959] = 92;
// bram[26960] = 76;
// bram[26961] = 61;
// bram[26962] = 46;
// bram[26963] = 34;
// bram[26964] = 23;
// bram[26965] = 14;
// bram[26966] = 7;
// bram[26967] = 2;
// bram[26968] = 0;
// bram[26969] = 0;
// bram[26970] = 2;
// bram[26971] = 7;
// bram[26972] = 14;
// bram[26973] = 23;
// bram[26974] = 34;
// bram[26975] = 47;
// bram[26976] = 61;
// bram[26977] = 77;
// bram[26978] = 93;
// bram[26979] = 110;
// bram[26980] = 127;
// bram[26981] = 145;
// bram[26982] = 162;
// bram[26983] = 178;
// bram[26984] = 194;
// bram[26985] = 208;
// bram[26986] = 220;
// bram[26987] = 231;
// bram[26988] = 240;
// bram[26989] = 247;
// bram[26990] = 251;
// bram[26991] = 253;
// bram[26992] = 253;
// bram[26993] = 250;
// bram[26994] = 246;
// bram[26995] = 238;
// bram[26996] = 229;
// bram[26997] = 218;
// bram[26998] = 205;
// bram[26999] = 191;
// bram[27000] = 175;
// bram[27001] = 159;
// bram[27002] = 142;
// bram[27003] = 124;
// bram[27004] = 107;
// bram[27005] = 90;
// bram[27006] = 74;
// bram[27007] = 58;
// bram[27008] = 44;
// bram[27009] = 32;
// bram[27010] = 21;
// bram[27011] = 12;
// bram[27012] = 6;
// bram[27013] = 2;
// bram[27014] = 0;
// bram[27015] = 0;
// bram[27016] = 3;
// bram[27017] = 8;
// bram[27018] = 15;
// bram[27019] = 25;
// bram[27020] = 36;
// bram[27021] = 49;
// bram[27022] = 63;
// bram[27023] = 79;
// bram[27024] = 96;
// bram[27025] = 113;
// bram[27026] = 130;
// bram[27027] = 147;
// bram[27028] = 164;
// bram[27029] = 181;
// bram[27030] = 196;
// bram[27031] = 210;
// bram[27032] = 222;
// bram[27033] = 233;
// bram[27034] = 241;
// bram[27035] = 248;
// bram[27036] = 252;
// bram[27037] = 253;
// bram[27038] = 253;
// bram[27039] = 250;
// bram[27040] = 245;
// bram[27041] = 237;
// bram[27042] = 228;
// bram[27043] = 216;
// bram[27044] = 203;
// bram[27045] = 188;
// bram[27046] = 173;
// bram[27047] = 156;
// bram[27048] = 139;
// bram[27049] = 121;
// bram[27050] = 104;
// bram[27051] = 87;
// bram[27052] = 71;
// bram[27053] = 56;
// bram[27054] = 42;
// bram[27055] = 30;
// bram[27056] = 20;
// bram[27057] = 11;
// bram[27058] = 5;
// bram[27059] = 1;
// bram[27060] = 0;
// bram[27061] = 0;
// bram[27062] = 3;
// bram[27063] = 9;
// bram[27064] = 17;
// bram[27065] = 26;
// bram[27066] = 38;
// bram[27067] = 51;
// bram[27068] = 66;
// bram[27069] = 82;
// bram[27070] = 98;
// bram[27071] = 115;
// bram[27072] = 133;
// bram[27073] = 150;
// bram[27074] = 167;
// bram[27075] = 183;
// bram[27076] = 198;
// bram[27077] = 212;
// bram[27078] = 224;
// bram[27079] = 234;
// bram[27080] = 242;
// bram[27081] = 248;
// bram[27082] = 252;
// bram[27083] = 253;
// bram[27084] = 253;
// bram[27085] = 249;
// bram[27086] = 244;
// bram[27087] = 236;
// bram[27088] = 226;
// bram[27089] = 214;
// bram[27090] = 201;
// bram[27091] = 186;
// bram[27092] = 170;
// bram[27093] = 153;
// bram[27094] = 136;
// bram[27095] = 119;
// bram[27096] = 102;
// bram[27097] = 85;
// bram[27098] = 69;
// bram[27099] = 54;
// bram[27100] = 40;
// bram[27101] = 28;
// bram[27102] = 18;
// bram[27103] = 10;
// bram[27104] = 4;
// bram[27105] = 1;
// bram[27106] = 0;
// bram[27107] = 1;
// bram[27108] = 4;
// bram[27109] = 10;
// bram[27110] = 18;
// bram[27111] = 28;
// bram[27112] = 40;
// bram[27113] = 53;
// bram[27114] = 68;
// bram[27115] = 84;
// bram[27116] = 101;
// bram[27117] = 118;
// bram[27118] = 136;
// bram[27119] = 153;
// bram[27120] = 170;
// bram[27121] = 185;
// bram[27122] = 200;
// bram[27123] = 214;
// bram[27124] = 225;
// bram[27125] = 235;
// bram[27126] = 243;
// bram[27127] = 249;
// bram[27128] = 252;
// bram[27129] = 253;
// bram[27130] = 252;
// bram[27131] = 248;
// bram[27132] = 242;
// bram[27133] = 234;
// bram[27134] = 224;
// bram[27135] = 212;
// bram[27136] = 199;
// bram[27137] = 184;
// bram[27138] = 168;
// bram[27139] = 151;
// bram[27140] = 133;
// bram[27141] = 116;
// bram[27142] = 99;
// bram[27143] = 82;
// bram[27144] = 66;
// bram[27145] = 52;
// bram[27146] = 38;
// bram[27147] = 27;
// bram[27148] = 17;
// bram[27149] = 9;
// bram[27150] = 4;
// bram[27151] = 0;
// bram[27152] = 0;
// bram[27153] = 1;
// bram[27154] = 5;
// bram[27155] = 11;
// bram[27156] = 19;
// bram[27157] = 30;
// bram[27158] = 42;
// bram[27159] = 56;
// bram[27160] = 71;
// bram[27161] = 87;
// bram[27162] = 104;
// bram[27163] = 121;
// bram[27164] = 138;
// bram[27165] = 155;
// bram[27166] = 172;
// bram[27167] = 188;
// bram[27168] = 202;
// bram[27169] = 216;
// bram[27170] = 227;
// bram[27171] = 237;
// bram[27172] = 244;
// bram[27173] = 250;
// bram[27174] = 253;
// bram[27175] = 253;
// bram[27176] = 252;
// bram[27177] = 248;
// bram[27178] = 241;
// bram[27179] = 233;
// bram[27180] = 222;
// bram[27181] = 210;
// bram[27182] = 196;
// bram[27183] = 181;
// bram[27184] = 165;
// bram[27185] = 148;
// bram[27186] = 131;
// bram[27187] = 113;
// bram[27188] = 96;
// bram[27189] = 80;
// bram[27190] = 64;
// bram[27191] = 49;
// bram[27192] = 36;
// bram[27193] = 25;
// bram[27194] = 16;
// bram[27195] = 8;
// bram[27196] = 3;
// bram[27197] = 0;
// bram[27198] = 0;
// bram[27199] = 1;
// bram[27200] = 6;
// bram[27201] = 12;
// bram[27202] = 21;
// bram[27203] = 31;
// bram[27204] = 44;
// bram[27205] = 58;
// bram[27206] = 73;
// bram[27207] = 89;
// bram[27208] = 106;
// bram[27209] = 124;
// bram[27210] = 141;
// bram[27211] = 158;
// bram[27212] = 175;
// bram[27213] = 190;
// bram[27214] = 205;
// bram[27215] = 218;
// bram[27216] = 229;
// bram[27217] = 238;
// bram[27218] = 245;
// bram[27219] = 250;
// bram[27220] = 253;
// bram[27221] = 253;
// bram[27222] = 251;
// bram[27223] = 247;
// bram[27224] = 240;
// bram[27225] = 231;
// bram[27226] = 221;
// bram[27227] = 208;
// bram[27228] = 194;
// bram[27229] = 179;
// bram[27230] = 162;
// bram[27231] = 145;
// bram[27232] = 128;
// bram[27233] = 111;
// bram[27234] = 94;
// bram[27235] = 77;
// bram[27236] = 62;
// bram[27237] = 47;
// bram[27238] = 35;
// bram[27239] = 23;
// bram[27240] = 14;
// bram[27241] = 7;
// bram[27242] = 2;
// bram[27243] = 0;
// bram[27244] = 0;
// bram[27245] = 2;
// bram[27246] = 7;
// bram[27247] = 13;
// bram[27248] = 22;
// bram[27249] = 33;
// bram[27250] = 46;
// bram[27251] = 60;
// bram[27252] = 76;
// bram[27253] = 92;
// bram[27254] = 109;
// bram[27255] = 126;
// bram[27256] = 144;
// bram[27257] = 161;
// bram[27258] = 177;
// bram[27259] = 192;
// bram[27260] = 207;
// bram[27261] = 219;
// bram[27262] = 230;
// bram[27263] = 239;
// bram[27264] = 246;
// bram[27265] = 251;
// bram[27266] = 253;
// bram[27267] = 253;
// bram[27268] = 251;
// bram[27269] = 246;
// bram[27270] = 239;
// bram[27271] = 230;
// bram[27272] = 219;
// bram[27273] = 206;
// bram[27274] = 192;
// bram[27275] = 176;
// bram[27276] = 160;
// bram[27277] = 143;
// bram[27278] = 125;
// bram[27279] = 108;
// bram[27280] = 91;
// bram[27281] = 75;
// bram[27282] = 59;
// bram[27283] = 45;
// bram[27284] = 33;
// bram[27285] = 22;
// bram[27286] = 13;
// bram[27287] = 6;
// bram[27288] = 2;
// bram[27289] = 0;
// bram[27290] = 0;
// bram[27291] = 3;
// bram[27292] = 7;
// bram[27293] = 15;
// bram[27294] = 24;
// bram[27295] = 35;
// bram[27296] = 48;
// bram[27297] = 62;
// bram[27298] = 78;
// bram[27299] = 94;
// bram[27300] = 112;
// bram[27301] = 129;
// bram[27302] = 146;
// bram[27303] = 163;
// bram[27304] = 179;
// bram[27305] = 195;
// bram[27306] = 209;
// bram[27307] = 221;
// bram[27308] = 232;
// bram[27309] = 241;
// bram[27310] = 247;
// bram[27311] = 251;
// bram[27312] = 253;
// bram[27313] = 253;
// bram[27314] = 250;
// bram[27315] = 245;
// bram[27316] = 238;
// bram[27317] = 228;
// bram[27318] = 217;
// bram[27319] = 204;
// bram[27320] = 189;
// bram[27321] = 174;
// bram[27322] = 157;
// bram[27323] = 140;
// bram[27324] = 123;
// bram[27325] = 105;
// bram[27326] = 88;
// bram[27327] = 72;
// bram[27328] = 57;
// bram[27329] = 43;
// bram[27330] = 31;
// bram[27331] = 20;
// bram[27332] = 12;
// bram[27333] = 5;
// bram[27334] = 1;
// bram[27335] = 0;
// bram[27336] = 0;
// bram[27337] = 3;
// bram[27338] = 8;
// bram[27339] = 16;
// bram[27340] = 26;
// bram[27341] = 37;
// bram[27342] = 50;
// bram[27343] = 65;
// bram[27344] = 80;
// bram[27345] = 97;
// bram[27346] = 114;
// bram[27347] = 132;
// bram[27348] = 149;
// bram[27349] = 166;
// bram[27350] = 182;
// bram[27351] = 197;
// bram[27352] = 211;
// bram[27353] = 223;
// bram[27354] = 233;
// bram[27355] = 242;
// bram[27356] = 248;
// bram[27357] = 252;
// bram[27358] = 253;
// bram[27359] = 253;
// bram[27360] = 250;
// bram[27361] = 244;
// bram[27362] = 236;
// bram[27363] = 227;
// bram[27364] = 215;
// bram[27365] = 202;
// bram[27366] = 187;
// bram[27367] = 171;
// bram[27368] = 155;
// bram[27369] = 137;
// bram[27370] = 120;
// bram[27371] = 103;
// bram[27372] = 86;
// bram[27373] = 70;
// bram[27374] = 55;
// bram[27375] = 41;
// bram[27376] = 29;
// bram[27377] = 19;
// bram[27378] = 11;
// bram[27379] = 5;
// bram[27380] = 1;
// bram[27381] = 0;
// bram[27382] = 0;
// bram[27383] = 4;
// bram[27384] = 9;
// bram[27385] = 17;
// bram[27386] = 27;
// bram[27387] = 39;
// bram[27388] = 52;
// bram[27389] = 67;
// bram[27390] = 83;
// bram[27391] = 100;
// bram[27392] = 117;
// bram[27393] = 134;
// bram[27394] = 152;
// bram[27395] = 168;
// bram[27396] = 184;
// bram[27397] = 199;
// bram[27398] = 213;
// bram[27399] = 225;
// bram[27400] = 235;
// bram[27401] = 243;
// bram[27402] = 249;
// bram[27403] = 252;
// bram[27404] = 253;
// bram[27405] = 252;
// bram[27406] = 249;
// bram[27407] = 243;
// bram[27408] = 235;
// bram[27409] = 225;
// bram[27410] = 213;
// bram[27411] = 200;
// bram[27412] = 185;
// bram[27413] = 169;
// bram[27414] = 152;
// bram[27415] = 135;
// bram[27416] = 117;
// bram[27417] = 100;
// bram[27418] = 83;
// bram[27419] = 67;
// bram[27420] = 53;
// bram[27421] = 39;
// bram[27422] = 27;
// bram[27423] = 18;
// bram[27424] = 10;
// bram[27425] = 4;
// bram[27426] = 1;
// bram[27427] = 0;
// bram[27428] = 1;
// bram[27429] = 5;
// bram[27430] = 11;
// bram[27431] = 19;
// bram[27432] = 29;
// bram[27433] = 41;
// bram[27434] = 55;
// bram[27435] = 70;
// bram[27436] = 86;
// bram[27437] = 102;
// bram[27438] = 120;
// bram[27439] = 137;
// bram[27440] = 154;
// bram[27441] = 171;
// bram[27442] = 187;
// bram[27443] = 201;
// bram[27444] = 215;
// bram[27445] = 226;
// bram[27446] = 236;
// bram[27447] = 244;
// bram[27448] = 249;
// bram[27449] = 253;
// bram[27450] = 253;
// bram[27451] = 252;
// bram[27452] = 248;
// bram[27453] = 242;
// bram[27454] = 234;
// bram[27455] = 223;
// bram[27456] = 211;
// bram[27457] = 197;
// bram[27458] = 182;
// bram[27459] = 166;
// bram[27460] = 149;
// bram[27461] = 132;
// bram[27462] = 115;
// bram[27463] = 97;
// bram[27464] = 81;
// bram[27465] = 65;
// bram[27466] = 50;
// bram[27467] = 37;
// bram[27468] = 26;
// bram[27469] = 16;
// bram[27470] = 9;
// bram[27471] = 3;
// bram[27472] = 0;
// bram[27473] = 0;
// bram[27474] = 1;
// bram[27475] = 5;
// bram[27476] = 12;
// bram[27477] = 20;
// bram[27478] = 31;
// bram[27479] = 43;
// bram[27480] = 57;
// bram[27481] = 72;
// bram[27482] = 88;
// bram[27483] = 105;
// bram[27484] = 122;
// bram[27485] = 140;
// bram[27486] = 157;
// bram[27487] = 173;
// bram[27488] = 189;
// bram[27489] = 204;
// bram[27490] = 217;
// bram[27491] = 228;
// bram[27492] = 238;
// bram[27493] = 245;
// bram[27494] = 250;
// bram[27495] = 253;
// bram[27496] = 253;
// bram[27497] = 251;
// bram[27498] = 247;
// bram[27499] = 241;
// bram[27500] = 232;
// bram[27501] = 221;
// bram[27502] = 209;
// bram[27503] = 195;
// bram[27504] = 180;
// bram[27505] = 164;
// bram[27506] = 147;
// bram[27507] = 129;
// bram[27508] = 112;
// bram[27509] = 95;
// bram[27510] = 78;
// bram[27511] = 63;
// bram[27512] = 48;
// bram[27513] = 35;
// bram[27514] = 24;
// bram[27515] = 15;
// bram[27516] = 8;
// bram[27517] = 3;
// bram[27518] = 0;
// bram[27519] = 0;
// bram[27520] = 2;
// bram[27521] = 6;
// bram[27522] = 13;
// bram[27523] = 22;
// bram[27524] = 32;
// bram[27525] = 45;
// bram[27526] = 59;
// bram[27527] = 74;
// bram[27528] = 91;
// bram[27529] = 108;
// bram[27530] = 125;
// bram[27531] = 142;
// bram[27532] = 159;
// bram[27533] = 176;
// bram[27534] = 191;
// bram[27535] = 206;
// bram[27536] = 219;
// bram[27537] = 230;
// bram[27538] = 239;
// bram[27539] = 246;
// bram[27540] = 251;
// bram[27541] = 253;
// bram[27542] = 253;
// bram[27543] = 251;
// bram[27544] = 246;
// bram[27545] = 240;
// bram[27546] = 231;
// bram[27547] = 220;
// bram[27548] = 207;
// bram[27549] = 193;
// bram[27550] = 177;
// bram[27551] = 161;
// bram[27552] = 144;
// bram[27553] = 127;
// bram[27554] = 109;
// bram[27555] = 92;
// bram[27556] = 76;
// bram[27557] = 60;
// bram[27558] = 46;
// bram[27559] = 34;
// bram[27560] = 23;
// bram[27561] = 14;
// bram[27562] = 7;
// bram[27563] = 2;
// bram[27564] = 0;
// bram[27565] = 0;
// bram[27566] = 2;
// bram[27567] = 7;
// bram[27568] = 14;
// bram[27569] = 23;
// bram[27570] = 34;
// bram[27571] = 47;
// bram[27572] = 61;
// bram[27573] = 77;
// bram[27574] = 93;
// bram[27575] = 110;
// bram[27576] = 128;
// bram[27577] = 145;
// bram[27578] = 162;
// bram[27579] = 178;
// bram[27580] = 194;
// bram[27581] = 208;
// bram[27582] = 220;
// bram[27583] = 231;
// bram[27584] = 240;
// bram[27585] = 247;
// bram[27586] = 251;
// bram[27587] = 253;
// bram[27588] = 253;
// bram[27589] = 250;
// bram[27590] = 245;
// bram[27591] = 238;
// bram[27592] = 229;
// bram[27593] = 218;
// bram[27594] = 205;
// bram[27595] = 191;
// bram[27596] = 175;
// bram[27597] = 158;
// bram[27598] = 141;
// bram[27599] = 124;
// bram[27600] = 107;
// bram[27601] = 90;
// bram[27602] = 73;
// bram[27603] = 58;
// bram[27604] = 44;
// bram[27605] = 32;
// bram[27606] = 21;
// bram[27607] = 12;
// bram[27608] = 6;
// bram[27609] = 2;
// bram[27610] = 0;
// bram[27611] = 0;
// bram[27612] = 3;
// bram[27613] = 8;
// bram[27614] = 15;
// bram[27615] = 25;
// bram[27616] = 36;
// bram[27617] = 49;
// bram[27618] = 64;
// bram[27619] = 79;
// bram[27620] = 96;
// bram[27621] = 113;
// bram[27622] = 130;
// bram[27623] = 148;
// bram[27624] = 165;
// bram[27625] = 181;
// bram[27626] = 196;
// bram[27627] = 210;
// bram[27628] = 222;
// bram[27629] = 233;
// bram[27630] = 241;
// bram[27631] = 248;
// bram[27632] = 252;
// bram[27633] = 253;
// bram[27634] = 253;
// bram[27635] = 250;
// bram[27636] = 245;
// bram[27637] = 237;
// bram[27638] = 227;
// bram[27639] = 216;
// bram[27640] = 203;
// bram[27641] = 188;
// bram[27642] = 172;
// bram[27643] = 156;
// bram[27644] = 139;
// bram[27645] = 121;
// bram[27646] = 104;
// bram[27647] = 87;
// bram[27648] = 71;
// bram[27649] = 56;
// bram[27650] = 42;
// bram[27651] = 30;
// bram[27652] = 20;
// bram[27653] = 11;
// bram[27654] = 5;
// bram[27655] = 1;
// bram[27656] = 0;
// bram[27657] = 0;
// bram[27658] = 4;
// bram[27659] = 9;
// bram[27660] = 17;
// bram[27661] = 26;
// bram[27662] = 38;
// bram[27663] = 51;
// bram[27664] = 66;
// bram[27665] = 82;
// bram[27666] = 99;
// bram[27667] = 116;
// bram[27668] = 133;
// bram[27669] = 150;
// bram[27670] = 167;
// bram[27671] = 183;
// bram[27672] = 198;
// bram[27673] = 212;
// bram[27674] = 224;
// bram[27675] = 234;
// bram[27676] = 242;
// bram[27677] = 248;
// bram[27678] = 252;
// bram[27679] = 253;
// bram[27680] = 252;
// bram[27681] = 249;
// bram[27682] = 243;
// bram[27683] = 236;
// bram[27684] = 226;
// bram[27685] = 214;
// bram[27686] = 201;
// bram[27687] = 186;
// bram[27688] = 170;
// bram[27689] = 153;
// bram[27690] = 136;
// bram[27691] = 119;
// bram[27692] = 101;
// bram[27693] = 85;
// bram[27694] = 69;
// bram[27695] = 54;
// bram[27696] = 40;
// bram[27697] = 28;
// bram[27698] = 18;
// bram[27699] = 10;
// bram[27700] = 4;
// bram[27701] = 1;
// bram[27702] = 0;
// bram[27703] = 1;
// bram[27704] = 4;
// bram[27705] = 10;
// bram[27706] = 18;
// bram[27707] = 28;
// bram[27708] = 40;
// bram[27709] = 54;
// bram[27710] = 68;
// bram[27711] = 84;
// bram[27712] = 101;
// bram[27713] = 118;
// bram[27714] = 136;
// bram[27715] = 153;
// bram[27716] = 170;
// bram[27717] = 186;
// bram[27718] = 200;
// bram[27719] = 214;
// bram[27720] = 226;
// bram[27721] = 236;
// bram[27722] = 243;
// bram[27723] = 249;
// bram[27724] = 252;
// bram[27725] = 253;
// bram[27726] = 252;
// bram[27727] = 248;
// bram[27728] = 242;
// bram[27729] = 234;
// bram[27730] = 224;
// bram[27731] = 212;
// bram[27732] = 198;
// bram[27733] = 183;
// bram[27734] = 167;
// bram[27735] = 151;
// bram[27736] = 133;
// bram[27737] = 116;
// bram[27738] = 99;
// bram[27739] = 82;
// bram[27740] = 66;
// bram[27741] = 51;
// bram[27742] = 38;
// bram[27743] = 27;
// bram[27744] = 17;
// bram[27745] = 9;
// bram[27746] = 4;
// bram[27747] = 0;
// bram[27748] = 0;
// bram[27749] = 1;
// bram[27750] = 5;
// bram[27751] = 11;
// bram[27752] = 19;
// bram[27753] = 30;
// bram[27754] = 42;
// bram[27755] = 56;
// bram[27756] = 71;
// bram[27757] = 87;
// bram[27758] = 104;
// bram[27759] = 121;
// bram[27760] = 138;
// bram[27761] = 156;
// bram[27762] = 172;
// bram[27763] = 188;
// bram[27764] = 203;
// bram[27765] = 216;
// bram[27766] = 227;
// bram[27767] = 237;
// bram[27768] = 244;
// bram[27769] = 250;
// bram[27770] = 253;
// bram[27771] = 253;
// bram[27772] = 252;
// bram[27773] = 248;
// bram[27774] = 241;
// bram[27775] = 233;
// bram[27776] = 222;
// bram[27777] = 210;
// bram[27778] = 196;
// bram[27779] = 181;
// bram[27780] = 165;
// bram[27781] = 148;
// bram[27782] = 131;
// bram[27783] = 113;
// bram[27784] = 96;
// bram[27785] = 80;
// bram[27786] = 64;
// bram[27787] = 49;
// bram[27788] = 36;
// bram[27789] = 25;
// bram[27790] = 15;
// bram[27791] = 8;
// bram[27792] = 3;
// bram[27793] = 0;
// bram[27794] = 0;
// bram[27795] = 2;
// bram[27796] = 6;
// bram[27797] = 12;
// bram[27798] = 21;
// bram[27799] = 32;
// bram[27800] = 44;
// bram[27801] = 58;
// bram[27802] = 73;
// bram[27803] = 89;
// bram[27804] = 106;
// bram[27805] = 124;
// bram[27806] = 141;
// bram[27807] = 158;
// bram[27808] = 175;
// bram[27809] = 190;
// bram[27810] = 205;
// bram[27811] = 218;
// bram[27812] = 229;
// bram[27813] = 238;
// bram[27814] = 245;
// bram[27815] = 250;
// bram[27816] = 253;
// bram[27817] = 253;
// bram[27818] = 251;
// bram[27819] = 247;
// bram[27820] = 240;
// bram[27821] = 231;
// bram[27822] = 221;
// bram[27823] = 208;
// bram[27824] = 194;
// bram[27825] = 179;
// bram[27826] = 162;
// bram[27827] = 145;
// bram[27828] = 128;
// bram[27829] = 111;
// bram[27830] = 93;
// bram[27831] = 77;
// bram[27832] = 62;
// bram[27833] = 47;
// bram[27834] = 34;
// bram[27835] = 23;
// bram[27836] = 14;
// bram[27837] = 7;
// bram[27838] = 2;
// bram[27839] = 0;
// bram[27840] = 0;
// bram[27841] = 2;
// bram[27842] = 7;
// bram[27843] = 14;
// bram[27844] = 22;
// bram[27845] = 33;
// bram[27846] = 46;
// bram[27847] = 60;
// bram[27848] = 76;
// bram[27849] = 92;
// bram[27850] = 109;
// bram[27851] = 126;
// bram[27852] = 144;
// bram[27853] = 161;
// bram[27854] = 177;
// bram[27855] = 193;
// bram[27856] = 207;
// bram[27857] = 220;
// bram[27858] = 230;
// bram[27859] = 239;
// bram[27860] = 246;
// bram[27861] = 251;
// bram[27862] = 253;
// bram[27863] = 253;
// bram[27864] = 251;
// bram[27865] = 246;
// bram[27866] = 239;
// bram[27867] = 230;
// bram[27868] = 219;
// bram[27869] = 206;
// bram[27870] = 192;
// bram[27871] = 176;
// bram[27872] = 160;
// bram[27873] = 143;
// bram[27874] = 125;
// bram[27875] = 108;
// bram[27876] = 91;
// bram[27877] = 75;
// bram[27878] = 59;
// bram[27879] = 45;
// bram[27880] = 33;
// bram[27881] = 22;
// bram[27882] = 13;
// bram[27883] = 6;
// bram[27884] = 2;
// bram[27885] = 0;
// bram[27886] = 0;
// bram[27887] = 3;
// bram[27888] = 8;
// bram[27889] = 15;
// bram[27890] = 24;
// bram[27891] = 35;
// bram[27892] = 48;
// bram[27893] = 63;
// bram[27894] = 78;
// bram[27895] = 95;
// bram[27896] = 112;
// bram[27897] = 129;
// bram[27898] = 146;
// bram[27899] = 163;
// bram[27900] = 180;
// bram[27901] = 195;
// bram[27902] = 209;
// bram[27903] = 221;
// bram[27904] = 232;
// bram[27905] = 241;
// bram[27906] = 247;
// bram[27907] = 251;
// bram[27908] = 253;
// bram[27909] = 253;
// bram[27910] = 250;
// bram[27911] = 245;
// bram[27912] = 238;
// bram[27913] = 228;
// bram[27914] = 217;
// bram[27915] = 204;
// bram[27916] = 189;
// bram[27917] = 174;
// bram[27918] = 157;
// bram[27919] = 140;
// bram[27920] = 123;
// bram[27921] = 105;
// bram[27922] = 88;
// bram[27923] = 72;
// bram[27924] = 57;
// bram[27925] = 43;
// bram[27926] = 31;
// bram[27927] = 20;
// bram[27928] = 12;
// bram[27929] = 5;
// bram[27930] = 1;
// bram[27931] = 0;
// bram[27932] = 0;
// bram[27933] = 3;
// bram[27934] = 9;
// bram[27935] = 16;
// bram[27936] = 26;
// bram[27937] = 37;
// bram[27938] = 50;
// bram[27939] = 65;
// bram[27940] = 81;
// bram[27941] = 97;
// bram[27942] = 114;
// bram[27943] = 132;
// bram[27944] = 149;
// bram[27945] = 166;
// bram[27946] = 182;
// bram[27947] = 197;
// bram[27948] = 211;
// bram[27949] = 223;
// bram[27950] = 233;
// bram[27951] = 242;
// bram[27952] = 248;
// bram[27953] = 252;
// bram[27954] = 253;
// bram[27955] = 253;
// bram[27956] = 249;
// bram[27957] = 244;
// bram[27958] = 236;
// bram[27959] = 227;
// bram[27960] = 215;
// bram[27961] = 202;
// bram[27962] = 187;
// bram[27963] = 171;
// bram[27964] = 154;
// bram[27965] = 137;
// bram[27966] = 120;
// bram[27967] = 103;
// bram[27968] = 86;
// bram[27969] = 70;
// bram[27970] = 55;
// bram[27971] = 41;
// bram[27972] = 29;
// bram[27973] = 19;
// bram[27974] = 11;
// bram[27975] = 5;
// bram[27976] = 1;
// bram[27977] = 0;
// bram[27978] = 1;
// bram[27979] = 4;
// bram[27980] = 10;
// bram[27981] = 17;
// bram[27982] = 27;
// bram[27983] = 39;
// bram[27984] = 52;
// bram[27985] = 67;
// bram[27986] = 83;
// bram[27987] = 100;
// bram[27988] = 117;
// bram[27989] = 135;
// bram[27990] = 152;
// bram[27991] = 169;
// bram[27992] = 185;
// bram[27993] = 199;
// bram[27994] = 213;
// bram[27995] = 225;
// bram[27996] = 235;
// bram[27997] = 243;
// bram[27998] = 249;
// bram[27999] = 252;
// bram[28000] = 254;
// bram[28001] = 252;
// bram[28002] = 249;
// bram[28003] = 243;
// bram[28004] = 235;
// bram[28005] = 225;
// bram[28006] = 213;
// bram[28007] = 199;
// bram[28008] = 185;
// bram[28009] = 169;
// bram[28010] = 152;
// bram[28011] = 135;
// bram[28012] = 117;
// bram[28013] = 100;
// bram[28014] = 83;
// bram[28015] = 67;
// bram[28016] = 52;
// bram[28017] = 39;
// bram[28018] = 27;
// bram[28019] = 17;
// bram[28020] = 10;
// bram[28021] = 4;
// bram[28022] = 1;
// bram[28023] = 0;
// bram[28024] = 1;
// bram[28025] = 5;
// bram[28026] = 11;
// bram[28027] = 19;
// bram[28028] = 29;
// bram[28029] = 41;
// bram[28030] = 55;
// bram[28031] = 70;
// bram[28032] = 86;
// bram[28033] = 103;
// bram[28034] = 120;
// bram[28035] = 137;
// bram[28036] = 154;
// bram[28037] = 171;
// bram[28038] = 187;
// bram[28039] = 202;
// bram[28040] = 215;
// bram[28041] = 227;
// bram[28042] = 236;
// bram[28043] = 244;
// bram[28044] = 249;
// bram[28045] = 253;
// bram[28046] = 253;
// bram[28047] = 252;
// bram[28048] = 248;
// bram[28049] = 242;
// bram[28050] = 233;
// bram[28051] = 223;
// bram[28052] = 211;
// bram[28053] = 197;
// bram[28054] = 182;
// bram[28055] = 166;
// bram[28056] = 149;
// bram[28057] = 132;
// bram[28058] = 114;
// bram[28059] = 97;
// bram[28060] = 81;
// bram[28061] = 65;
// bram[28062] = 50;
// bram[28063] = 37;
// bram[28064] = 26;
// bram[28065] = 16;
// bram[28066] = 9;
// bram[28067] = 3;
// bram[28068] = 0;
// bram[28069] = 0;
// bram[28070] = 1;
// bram[28071] = 5;
// bram[28072] = 12;
// bram[28073] = 20;
// bram[28074] = 31;
// bram[28075] = 43;
// bram[28076] = 57;
// bram[28077] = 72;
// bram[28078] = 88;
// bram[28079] = 105;
// bram[28080] = 123;
// bram[28081] = 140;
// bram[28082] = 157;
// bram[28083] = 174;
// bram[28084] = 189;
// bram[28085] = 204;
// bram[28086] = 217;
// bram[28087] = 228;
// bram[28088] = 238;
// bram[28089] = 245;
// bram[28090] = 250;
// bram[28091] = 253;
// bram[28092] = 253;
// bram[28093] = 251;
// bram[28094] = 247;
// bram[28095] = 241;
// bram[28096] = 232;
// bram[28097] = 221;
// bram[28098] = 209;
// bram[28099] = 195;
// bram[28100] = 180;
// bram[28101] = 163;
// bram[28102] = 146;
// bram[28103] = 129;
// bram[28104] = 112;
// bram[28105] = 95;
// bram[28106] = 78;
// bram[28107] = 63;
// bram[28108] = 48;
// bram[28109] = 35;
// bram[28110] = 24;
// bram[28111] = 15;
// bram[28112] = 8;
// bram[28113] = 3;
// bram[28114] = 0;
// bram[28115] = 0;
// bram[28116] = 2;
// bram[28117] = 6;
// bram[28118] = 13;
// bram[28119] = 22;
// bram[28120] = 33;
// bram[28121] = 45;
// bram[28122] = 59;
// bram[28123] = 75;
// bram[28124] = 91;
// bram[28125] = 108;
// bram[28126] = 125;
// bram[28127] = 143;
// bram[28128] = 160;
// bram[28129] = 176;
// bram[28130] = 192;
// bram[28131] = 206;
// bram[28132] = 219;
// bram[28133] = 230;
// bram[28134] = 239;
// bram[28135] = 246;
// bram[28136] = 251;
// bram[28137] = 253;
// bram[28138] = 253;
// bram[28139] = 251;
// bram[28140] = 246;
// bram[28141] = 239;
// bram[28142] = 230;
// bram[28143] = 220;
// bram[28144] = 207;
// bram[28145] = 193;
// bram[28146] = 177;
// bram[28147] = 161;
// bram[28148] = 144;
// bram[28149] = 126;
// bram[28150] = 109;
// bram[28151] = 92;
// bram[28152] = 76;
// bram[28153] = 60;
// bram[28154] = 46;
// bram[28155] = 33;
// bram[28156] = 22;
// bram[28157] = 14;
// bram[28158] = 7;
// bram[28159] = 2;
// bram[28160] = 0;
// bram[28161] = 0;
// bram[28162] = 2;
// bram[28163] = 7;
// bram[28164] = 14;
// bram[28165] = 23;
// bram[28166] = 34;
// bram[28167] = 47;
// bram[28168] = 62;
// bram[28169] = 77;
// bram[28170] = 93;
// bram[28171] = 111;
// bram[28172] = 128;
// bram[28173] = 145;
// bram[28174] = 162;
// bram[28175] = 179;
// bram[28176] = 194;
// bram[28177] = 208;
// bram[28178] = 221;
// bram[28179] = 231;
// bram[28180] = 240;
// bram[28181] = 247;
// bram[28182] = 251;
// bram[28183] = 253;
// bram[28184] = 253;
// bram[28185] = 250;
// bram[28186] = 245;
// bram[28187] = 238;
// bram[28188] = 229;
// bram[28189] = 218;
// bram[28190] = 205;
// bram[28191] = 190;
// bram[28192] = 175;
// bram[28193] = 158;
// bram[28194] = 141;
// bram[28195] = 124;
// bram[28196] = 106;
// bram[28197] = 89;
// bram[28198] = 73;
// bram[28199] = 58;
// bram[28200] = 44;
// bram[28201] = 32;
// bram[28202] = 21;
// bram[28203] = 12;
// bram[28204] = 6;
// bram[28205] = 2;
// bram[28206] = 0;
// bram[28207] = 0;
// bram[28208] = 3;
// bram[28209] = 8;
// bram[28210] = 15;
// bram[28211] = 25;
// bram[28212] = 36;
// bram[28213] = 49;
// bram[28214] = 64;
// bram[28215] = 80;
// bram[28216] = 96;
// bram[28217] = 113;
// bram[28218] = 131;
// bram[28219] = 148;
// bram[28220] = 165;
// bram[28221] = 181;
// bram[28222] = 196;
// bram[28223] = 210;
// bram[28224] = 222;
// bram[28225] = 233;
// bram[28226] = 241;
// bram[28227] = 248;
// bram[28228] = 252;
// bram[28229] = 253;
// bram[28230] = 253;
// bram[28231] = 250;
// bram[28232] = 244;
// bram[28233] = 237;
// bram[28234] = 227;
// bram[28235] = 216;
// bram[28236] = 203;
// bram[28237] = 188;
// bram[28238] = 172;
// bram[28239] = 156;
// bram[28240] = 138;
// bram[28241] = 121;
// bram[28242] = 104;
// bram[28243] = 87;
// bram[28244] = 71;
// bram[28245] = 56;
// bram[28246] = 42;
// bram[28247] = 30;
// bram[28248] = 19;
// bram[28249] = 11;
// bram[28250] = 5;
// bram[28251] = 1;
// bram[28252] = 0;
// bram[28253] = 0;
// bram[28254] = 4;
// bram[28255] = 9;
// bram[28256] = 17;
// bram[28257] = 27;
// bram[28258] = 38;
// bram[28259] = 51;
// bram[28260] = 66;
// bram[28261] = 82;
// bram[28262] = 99;
// bram[28263] = 116;
// bram[28264] = 133;
// bram[28265] = 151;
// bram[28266] = 167;
// bram[28267] = 183;
// bram[28268] = 198;
// bram[28269] = 212;
// bram[28270] = 224;
// bram[28271] = 234;
// bram[28272] = 242;
// bram[28273] = 248;
// bram[28274] = 252;
// bram[28275] = 253;
// bram[28276] = 252;
// bram[28277] = 249;
// bram[28278] = 243;
// bram[28279] = 236;
// bram[28280] = 226;
// bram[28281] = 214;
// bram[28282] = 200;
// bram[28283] = 186;
// bram[28284] = 170;
// bram[28285] = 153;
// bram[28286] = 136;
// bram[28287] = 118;
// bram[28288] = 101;
// bram[28289] = 84;
// bram[28290] = 68;
// bram[28291] = 54;
// bram[28292] = 40;
// bram[28293] = 28;
// bram[28294] = 18;
// bram[28295] = 10;
// bram[28296] = 4;
// bram[28297] = 1;
// bram[28298] = 0;
// bram[28299] = 1;
// bram[28300] = 4;
// bram[28301] = 10;
// bram[28302] = 18;
// bram[28303] = 28;
// bram[28304] = 40;
// bram[28305] = 54;
// bram[28306] = 69;
// bram[28307] = 85;
// bram[28308] = 101;
// bram[28309] = 119;
// bram[28310] = 136;
// bram[28311] = 153;
// bram[28312] = 170;
// bram[28313] = 186;
// bram[28314] = 201;
// bram[28315] = 214;
// bram[28316] = 226;
// bram[28317] = 236;
// bram[28318] = 243;
// bram[28319] = 249;
// bram[28320] = 252;
// bram[28321] = 253;
// bram[28322] = 252;
// bram[28323] = 248;
// bram[28324] = 242;
// bram[28325] = 234;
// bram[28326] = 224;
// bram[28327] = 212;
// bram[28328] = 198;
// bram[28329] = 183;
// bram[28330] = 167;
// bram[28331] = 150;
// bram[28332] = 133;
// bram[28333] = 116;
// bram[28334] = 99;
// bram[28335] = 82;
// bram[28336] = 66;
// bram[28337] = 51;
// bram[28338] = 38;
// bram[28339] = 26;
// bram[28340] = 17;
// bram[28341] = 9;
// bram[28342] = 4;
// bram[28343] = 0;
// bram[28344] = 0;
// bram[28345] = 1;
// bram[28346] = 5;
// bram[28347] = 11;
// bram[28348] = 20;
// bram[28349] = 30;
// bram[28350] = 42;
// bram[28351] = 56;
// bram[28352] = 71;
// bram[28353] = 87;
// bram[28354] = 104;
// bram[28355] = 121;
// bram[28356] = 139;
// bram[28357] = 156;
// bram[28358] = 172;
// bram[28359] = 188;
// bram[28360] = 203;
// bram[28361] = 216;
// bram[28362] = 227;
// bram[28363] = 237;
// bram[28364] = 245;
// bram[28365] = 250;
// bram[28366] = 253;
// bram[28367] = 253;
// bram[28368] = 252;
// bram[28369] = 248;
// bram[28370] = 241;
// bram[28371] = 233;
// bram[28372] = 222;
// bram[28373] = 210;
// bram[28374] = 196;
// bram[28375] = 181;
// bram[28376] = 165;
// bram[28377] = 148;
// bram[28378] = 130;
// bram[28379] = 113;
// bram[28380] = 96;
// bram[28381] = 79;
// bram[28382] = 64;
// bram[28383] = 49;
// bram[28384] = 36;
// bram[28385] = 25;
// bram[28386] = 15;
// bram[28387] = 8;
// bram[28388] = 3;
// bram[28389] = 0;
// bram[28390] = 0;
// bram[28391] = 2;
// bram[28392] = 6;
// bram[28393] = 12;
// bram[28394] = 21;
// bram[28395] = 32;
// bram[28396] = 44;
// bram[28397] = 58;
// bram[28398] = 73;
// bram[28399] = 90;
// bram[28400] = 107;
// bram[28401] = 124;
// bram[28402] = 141;
// bram[28403] = 158;
// bram[28404] = 175;
// bram[28405] = 191;
// bram[28406] = 205;
// bram[28407] = 218;
// bram[28408] = 229;
// bram[28409] = 238;
// bram[28410] = 245;
// bram[28411] = 250;
// bram[28412] = 253;
// bram[28413] = 253;
// bram[28414] = 251;
// bram[28415] = 247;
// bram[28416] = 240;
// bram[28417] = 231;
// bram[28418] = 220;
// bram[28419] = 208;
// bram[28420] = 194;
// bram[28421] = 178;
// bram[28422] = 162;
// bram[28423] = 145;
// bram[28424] = 128;
// bram[28425] = 110;
// bram[28426] = 93;
// bram[28427] = 77;
// bram[28428] = 61;
// bram[28429] = 47;
// bram[28430] = 34;
// bram[28431] = 23;
// bram[28432] = 14;
// bram[28433] = 7;
// bram[28434] = 2;
// bram[28435] = 0;
// bram[28436] = 0;
// bram[28437] = 2;
// bram[28438] = 7;
// bram[28439] = 14;
// bram[28440] = 23;
// bram[28441] = 34;
// bram[28442] = 46;
// bram[28443] = 60;
// bram[28444] = 76;
// bram[28445] = 92;
// bram[28446] = 109;
// bram[28447] = 127;
// bram[28448] = 144;
// bram[28449] = 161;
// bram[28450] = 177;
// bram[28451] = 193;
// bram[28452] = 207;
// bram[28453] = 220;
// bram[28454] = 231;
// bram[28455] = 240;
// bram[28456] = 246;
// bram[28457] = 251;
// bram[28458] = 253;
// bram[28459] = 253;
// bram[28460] = 251;
// bram[28461] = 246;
// bram[28462] = 239;
// bram[28463] = 230;
// bram[28464] = 219;
// bram[28465] = 206;
// bram[28466] = 191;
// bram[28467] = 176;
// bram[28468] = 159;
// bram[28469] = 142;
// bram[28470] = 125;
// bram[28471] = 108;
// bram[28472] = 91;
// bram[28473] = 74;
// bram[28474] = 59;
// bram[28475] = 45;
// bram[28476] = 32;
// bram[28477] = 22;
// bram[28478] = 13;
// bram[28479] = 6;
// bram[28480] = 2;
// bram[28481] = 0;
// bram[28482] = 0;
// bram[28483] = 3;
// bram[28484] = 8;
// bram[28485] = 15;
// bram[28486] = 24;
// bram[28487] = 35;
// bram[28488] = 48;
// bram[28489] = 63;
// bram[28490] = 78;
// bram[28491] = 95;
// bram[28492] = 112;
// bram[28493] = 129;
// bram[28494] = 147;
// bram[28495] = 164;
// bram[28496] = 180;
// bram[28497] = 195;
// bram[28498] = 209;
// bram[28499] = 221;
// bram[28500] = 232;
// bram[28501] = 241;
// bram[28502] = 247;
// bram[28503] = 251;
// bram[28504] = 253;
// bram[28505] = 253;
// bram[28506] = 250;
// bram[28507] = 245;
// bram[28508] = 238;
// bram[28509] = 228;
// bram[28510] = 217;
// bram[28511] = 204;
// bram[28512] = 189;
// bram[28513] = 173;
// bram[28514] = 157;
// bram[28515] = 140;
// bram[28516] = 122;
// bram[28517] = 105;
// bram[28518] = 88;
// bram[28519] = 72;
// bram[28520] = 57;
// bram[28521] = 43;
// bram[28522] = 31;
// bram[28523] = 20;
// bram[28524] = 12;
// bram[28525] = 5;
// bram[28526] = 1;
// bram[28527] = 0;
// bram[28528] = 0;
// bram[28529] = 3;
// bram[28530] = 9;
// bram[28531] = 16;
// bram[28532] = 26;
// bram[28533] = 37;
// bram[28534] = 50;
// bram[28535] = 65;
// bram[28536] = 81;
// bram[28537] = 97;
// bram[28538] = 115;
// bram[28539] = 132;
// bram[28540] = 149;
// bram[28541] = 166;
// bram[28542] = 182;
// bram[28543] = 197;
// bram[28544] = 211;
// bram[28545] = 223;
// bram[28546] = 234;
// bram[28547] = 242;
// bram[28548] = 248;
// bram[28549] = 252;
// bram[28550] = 253;
// bram[28551] = 253;
// bram[28552] = 249;
// bram[28553] = 244;
// bram[28554] = 236;
// bram[28555] = 226;
// bram[28556] = 215;
// bram[28557] = 201;
// bram[28558] = 187;
// bram[28559] = 171;
// bram[28560] = 154;
// bram[28561] = 137;
// bram[28562] = 120;
// bram[28563] = 102;
// bram[28564] = 86;
// bram[28565] = 70;
// bram[28566] = 55;
// bram[28567] = 41;
// bram[28568] = 29;
// bram[28569] = 19;
// bram[28570] = 11;
// bram[28571] = 5;
// bram[28572] = 1;
// bram[28573] = 0;
// bram[28574] = 1;
// bram[28575] = 4;
// bram[28576] = 10;
// bram[28577] = 18;
// bram[28578] = 27;
// bram[28579] = 39;
// bram[28580] = 53;
// bram[28581] = 67;
// bram[28582] = 83;
// bram[28583] = 100;
// bram[28584] = 117;
// bram[28585] = 135;
// bram[28586] = 152;
// bram[28587] = 169;
// bram[28588] = 185;
// bram[28589] = 200;
// bram[28590] = 213;
// bram[28591] = 225;
// bram[28592] = 235;
// bram[28593] = 243;
// bram[28594] = 249;
// bram[28595] = 252;
// bram[28596] = 253;
// bram[28597] = 252;
// bram[28598] = 249;
// bram[28599] = 243;
// bram[28600] = 235;
// bram[28601] = 225;
// bram[28602] = 213;
// bram[28603] = 199;
// bram[28604] = 184;
// bram[28605] = 168;
// bram[28606] = 152;
// bram[28607] = 134;
// bram[28608] = 117;
// bram[28609] = 100;
// bram[28610] = 83;
// bram[28611] = 67;
// bram[28612] = 52;
// bram[28613] = 39;
// bram[28614] = 27;
// bram[28615] = 17;
// bram[28616] = 9;
// bram[28617] = 4;
// bram[28618] = 0;
// bram[28619] = 0;
// bram[28620] = 1;
// bram[28621] = 5;
// bram[28622] = 11;
// bram[28623] = 19;
// bram[28624] = 29;
// bram[28625] = 41;
// bram[28626] = 55;
// bram[28627] = 70;
// bram[28628] = 86;
// bram[28629] = 103;
// bram[28630] = 120;
// bram[28631] = 137;
// bram[28632] = 155;
// bram[28633] = 171;
// bram[28634] = 187;
// bram[28635] = 202;
// bram[28636] = 215;
// bram[28637] = 227;
// bram[28638] = 236;
// bram[28639] = 244;
// bram[28640] = 250;
// bram[28641] = 253;
// bram[28642] = 253;
// bram[28643] = 252;
// bram[28644] = 248;
// bram[28645] = 242;
// bram[28646] = 233;
// bram[28647] = 223;
// bram[28648] = 211;
// bram[28649] = 197;
// bram[28650] = 182;
// bram[28651] = 166;
// bram[28652] = 149;
// bram[28653] = 132;
// bram[28654] = 114;
// bram[28655] = 97;
// bram[28656] = 80;
// bram[28657] = 65;
// bram[28658] = 50;
// bram[28659] = 37;
// bram[28660] = 26;
// bram[28661] = 16;
// bram[28662] = 8;
// bram[28663] = 3;
// bram[28664] = 0;
// bram[28665] = 0;
// bram[28666] = 1;
// bram[28667] = 5;
// bram[28668] = 12;
// bram[28669] = 20;
// bram[28670] = 31;
// bram[28671] = 43;
// bram[28672] = 57;
// bram[28673] = 72;
// bram[28674] = 88;
// bram[28675] = 105;
// bram[28676] = 123;
// bram[28677] = 140;
// bram[28678] = 157;
// bram[28679] = 174;
// bram[28680] = 189;
// bram[28681] = 204;
// bram[28682] = 217;
// bram[28683] = 228;
// bram[28684] = 238;
// bram[28685] = 245;
// bram[28686] = 250;
// bram[28687] = 253;
// bram[28688] = 253;
// bram[28689] = 251;
// bram[28690] = 247;
// bram[28691] = 241;
// bram[28692] = 232;
// bram[28693] = 221;
// bram[28694] = 209;
// bram[28695] = 195;
// bram[28696] = 179;
// bram[28697] = 163;
// bram[28698] = 146;
// bram[28699] = 129;
// bram[28700] = 112;
// bram[28701] = 94;
// bram[28702] = 78;
// bram[28703] = 62;
// bram[28704] = 48;
// bram[28705] = 35;
// bram[28706] = 24;
// bram[28707] = 15;
// bram[28708] = 7;
// bram[28709] = 3;
// bram[28710] = 0;
// bram[28711] = 0;
// bram[28712] = 2;
// bram[28713] = 6;
// bram[28714] = 13;
// bram[28715] = 22;
// bram[28716] = 33;
// bram[28717] = 45;
// bram[28718] = 59;
// bram[28719] = 75;
// bram[28720] = 91;
// bram[28721] = 108;
// bram[28722] = 125;
// bram[28723] = 143;
// bram[28724] = 160;
// bram[28725] = 176;
// bram[28726] = 192;
// bram[28727] = 206;
// bram[28728] = 219;
// bram[28729] = 230;
// bram[28730] = 239;
// bram[28731] = 246;
// bram[28732] = 251;
// bram[28733] = 253;
// bram[28734] = 253;
// bram[28735] = 251;
// bram[28736] = 246;
// bram[28737] = 239;
// bram[28738] = 230;
// bram[28739] = 219;
// bram[28740] = 207;
// bram[28741] = 192;
// bram[28742] = 177;
// bram[28743] = 161;
// bram[28744] = 144;
// bram[28745] = 126;
// bram[28746] = 109;
// bram[28747] = 92;
// bram[28748] = 76;
// bram[28749] = 60;
// bram[28750] = 46;
// bram[28751] = 33;
// bram[28752] = 22;
// bram[28753] = 13;
// bram[28754] = 7;
// bram[28755] = 2;
// bram[28756] = 0;
// bram[28757] = 0;
// bram[28758] = 2;
// bram[28759] = 7;
// bram[28760] = 14;
// bram[28761] = 23;
// bram[28762] = 35;
// bram[28763] = 47;
// bram[28764] = 62;
// bram[28765] = 77;
// bram[28766] = 94;
// bram[28767] = 111;
// bram[28768] = 128;
// bram[28769] = 145;
// bram[28770] = 162;
// bram[28771] = 179;
// bram[28772] = 194;
// bram[28773] = 208;
// bram[28774] = 221;
// bram[28775] = 231;
// bram[28776] = 240;
// bram[28777] = 247;
// bram[28778] = 251;
// bram[28779] = 253;
// bram[28780] = 253;
// bram[28781] = 250;
// bram[28782] = 245;
// bram[28783] = 238;
// bram[28784] = 229;
// bram[28785] = 218;
// bram[28786] = 205;
// bram[28787] = 190;
// bram[28788] = 175;
// bram[28789] = 158;
// bram[28790] = 141;
// bram[28791] = 124;
// bram[28792] = 106;
// bram[28793] = 89;
// bram[28794] = 73;
// bram[28795] = 58;
// bram[28796] = 44;
// bram[28797] = 31;
// bram[28798] = 21;
// bram[28799] = 12;
// bram[28800] = 6;
// bram[28801] = 1;
// bram[28802] = 0;
// bram[28803] = 0;
// bram[28804] = 3;
// bram[28805] = 8;
// bram[28806] = 16;
// bram[28807] = 25;
// bram[28808] = 36;
// bram[28809] = 49;
// bram[28810] = 64;
// bram[28811] = 80;
// bram[28812] = 96;
// bram[28813] = 113;
// bram[28814] = 131;
// bram[28815] = 148;
// bram[28816] = 165;
// bram[28817] = 181;
// bram[28818] = 196;
// bram[28819] = 210;
// bram[28820] = 222;
// bram[28821] = 233;
// bram[28822] = 241;
// bram[28823] = 248;
// bram[28824] = 252;
// bram[28825] = 253;
// bram[28826] = 253;
// bram[28827] = 250;
// bram[28828] = 244;
// bram[28829] = 237;
// bram[28830] = 227;
// bram[28831] = 216;
// bram[28832] = 202;
// bram[28833] = 188;
// bram[28834] = 172;
// bram[28835] = 155;
// bram[28836] = 138;
// bram[28837] = 121;
// bram[28838] = 104;
// bram[28839] = 87;
// bram[28840] = 71;
// bram[28841] = 56;
// bram[28842] = 42;
// bram[28843] = 30;
// bram[28844] = 19;
// bram[28845] = 11;
// bram[28846] = 5;
// bram[28847] = 1;
// bram[28848] = 0;
// bram[28849] = 0;
// bram[28850] = 4;
// bram[28851] = 9;
// bram[28852] = 17;
// bram[28853] = 27;
// bram[28854] = 38;
// bram[28855] = 52;
// bram[28856] = 66;
// bram[28857] = 82;
// bram[28858] = 99;
// bram[28859] = 116;
// bram[28860] = 133;
// bram[28861] = 151;
// bram[28862] = 168;
// bram[28863] = 184;
// bram[28864] = 199;
// bram[28865] = 212;
// bram[28866] = 224;
// bram[28867] = 234;
// bram[28868] = 242;
// bram[28869] = 248;
// bram[28870] = 252;
// bram[28871] = 253;
// bram[28872] = 252;
// bram[28873] = 249;
// bram[28874] = 243;
// bram[28875] = 235;
// bram[28876] = 225;
// bram[28877] = 214;
// bram[28878] = 200;
// bram[28879] = 185;
// bram[28880] = 170;
// bram[28881] = 153;
// bram[28882] = 136;
// bram[28883] = 118;
// bram[28884] = 101;
// bram[28885] = 84;
// bram[28886] = 68;
// bram[28887] = 53;
// bram[28888] = 40;
// bram[28889] = 28;
// bram[28890] = 18;
// bram[28891] = 10;
// bram[28892] = 4;
// bram[28893] = 1;
// bram[28894] = 0;
// bram[28895] = 1;
// bram[28896] = 4;
// bram[28897] = 10;
// bram[28898] = 18;
// bram[28899] = 28;
// bram[28900] = 40;
// bram[28901] = 54;
// bram[28902] = 69;
// bram[28903] = 85;
// bram[28904] = 102;
// bram[28905] = 119;
// bram[28906] = 136;
// bram[28907] = 153;
// bram[28908] = 170;
// bram[28909] = 186;
// bram[28910] = 201;
// bram[28911] = 214;
// bram[28912] = 226;
// bram[28913] = 236;
// bram[28914] = 244;
// bram[28915] = 249;
// bram[28916] = 253;
// bram[28917] = 253;
// bram[28918] = 252;
// bram[28919] = 248;
// bram[28920] = 242;
// bram[28921] = 234;
// bram[28922] = 224;
// bram[28923] = 212;
// bram[28924] = 198;
// bram[28925] = 183;
// bram[28926] = 167;
// bram[28927] = 150;
// bram[28928] = 133;
// bram[28929] = 115;
// bram[28930] = 98;
// bram[28931] = 82;
// bram[28932] = 66;
// bram[28933] = 51;
// bram[28934] = 38;
// bram[28935] = 26;
// bram[28936] = 17;
// bram[28937] = 9;
// bram[28938] = 3;
// bram[28939] = 0;
// bram[28940] = 0;
// bram[28941] = 1;
// bram[28942] = 5;
// bram[28943] = 11;
// bram[28944] = 20;
// bram[28945] = 30;
// bram[28946] = 42;
// bram[28947] = 56;
// bram[28948] = 71;
// bram[28949] = 87;
// bram[28950] = 104;
// bram[28951] = 121;
// bram[28952] = 139;
// bram[28953] = 156;
// bram[28954] = 173;
// bram[28955] = 188;
// bram[28956] = 203;
// bram[28957] = 216;
// bram[28958] = 228;
// bram[28959] = 237;
// bram[28960] = 245;
// bram[28961] = 250;
// bram[28962] = 253;
// bram[28963] = 253;
// bram[28964] = 252;
// bram[28965] = 248;
// bram[28966] = 241;
// bram[28967] = 233;
// bram[28968] = 222;
// bram[28969] = 210;
// bram[28970] = 196;
// bram[28971] = 181;
// bram[28972] = 164;
// bram[28973] = 147;
// bram[28974] = 130;
// bram[28975] = 113;
// bram[28976] = 96;
// bram[28977] = 79;
// bram[28978] = 63;
// bram[28979] = 49;
// bram[28980] = 36;
// bram[28981] = 25;
// bram[28982] = 15;
// bram[28983] = 8;
// bram[28984] = 3;
// bram[28985] = 0;
// bram[28986] = 0;
// bram[28987] = 2;
// bram[28988] = 6;
// bram[28989] = 12;
// bram[28990] = 21;
// bram[28991] = 32;
// bram[28992] = 44;
// bram[28993] = 58;
// bram[28994] = 74;
// bram[28995] = 90;
// bram[28996] = 107;
// bram[28997] = 124;
// bram[28998] = 142;
// bram[28999] = 159;
// bram[29000] = 175;
// bram[29001] = 191;
// bram[29002] = 205;
// bram[29003] = 218;
// bram[29004] = 229;
// bram[29005] = 238;
// bram[29006] = 246;
// bram[29007] = 250;
// bram[29008] = 253;
// bram[29009] = 253;
// bram[29010] = 251;
// bram[29011] = 247;
// bram[29012] = 240;
// bram[29013] = 231;
// bram[29014] = 220;
// bram[29015] = 208;
// bram[29016] = 194;
// bram[29017] = 178;
// bram[29018] = 162;
// bram[29019] = 145;
// bram[29020] = 127;
// bram[29021] = 110;
// bram[29022] = 93;
// bram[29023] = 77;
// bram[29024] = 61;
// bram[29025] = 47;
// bram[29026] = 34;
// bram[29027] = 23;
// bram[29028] = 14;
// bram[29029] = 7;
// bram[29030] = 2;
// bram[29031] = 0;
// bram[29032] = 0;
// bram[29033] = 2;
// bram[29034] = 7;
// bram[29035] = 14;
// bram[29036] = 23;
// bram[29037] = 34;
// bram[29038] = 46;
// bram[29039] = 61;
// bram[29040] = 76;
// bram[29041] = 92;
// bram[29042] = 109;
// bram[29043] = 127;
// bram[29044] = 144;
// bram[29045] = 161;
// bram[29046] = 178;
// bram[29047] = 193;
// bram[29048] = 207;
// bram[29049] = 220;
// bram[29050] = 231;
// bram[29051] = 240;
// bram[29052] = 246;
// bram[29053] = 251;
// bram[29054] = 253;
// bram[29055] = 253;
// bram[29056] = 251;
// bram[29057] = 246;
// bram[29058] = 239;
// bram[29059] = 230;
// bram[29060] = 218;
// bram[29061] = 206;
// bram[29062] = 191;
// bram[29063] = 176;
// bram[29064] = 159;
// bram[29065] = 142;
// bram[29066] = 125;
// bram[29067] = 107;
// bram[29068] = 90;
// bram[29069] = 74;
// bram[29070] = 59;
// bram[29071] = 45;
// bram[29072] = 32;
// bram[29073] = 22;
// bram[29074] = 13;
// bram[29075] = 6;
// bram[29076] = 2;
// bram[29077] = 0;
// bram[29078] = 0;
// bram[29079] = 3;
// bram[29080] = 8;
// bram[29081] = 15;
// bram[29082] = 24;
// bram[29083] = 36;
// bram[29084] = 49;
// bram[29085] = 63;
// bram[29086] = 79;
// bram[29087] = 95;
// bram[29088] = 112;
// bram[29089] = 130;
// bram[29090] = 147;
// bram[29091] = 164;
// bram[29092] = 180;
// bram[29093] = 195;
// bram[29094] = 209;
// bram[29095] = 222;
// bram[29096] = 232;
// bram[29097] = 241;
// bram[29098] = 247;
// bram[29099] = 252;
// bram[29100] = 253;
// bram[29101] = 253;
// bram[29102] = 250;
// bram[29103] = 245;
// bram[29104] = 237;
// bram[29105] = 228;
// bram[29106] = 217;
// bram[29107] = 203;
// bram[29108] = 189;
// bram[29109] = 173;
// bram[29110] = 157;
// bram[29111] = 139;
// bram[29112] = 122;
// bram[29113] = 105;
// bram[29114] = 88;
// bram[29115] = 72;
// bram[29116] = 57;
// bram[29117] = 43;
// bram[29118] = 31;
// bram[29119] = 20;
// bram[29120] = 12;
// bram[29121] = 5;
// bram[29122] = 1;
// bram[29123] = 0;
// bram[29124] = 0;
// bram[29125] = 3;
// bram[29126] = 9;
// bram[29127] = 16;
// bram[29128] = 26;
// bram[29129] = 37;
// bram[29130] = 51;
// bram[29131] = 65;
// bram[29132] = 81;
// bram[29133] = 98;
// bram[29134] = 115;
// bram[29135] = 132;
// bram[29136] = 150;
// bram[29137] = 166;
// bram[29138] = 182;
// bram[29139] = 198;
// bram[29140] = 211;
// bram[29141] = 223;
// bram[29142] = 234;
// bram[29143] = 242;
// bram[29144] = 248;
// bram[29145] = 252;
// bram[29146] = 253;
// bram[29147] = 253;
// bram[29148] = 249;
// bram[29149] = 244;
// bram[29150] = 236;
// bram[29151] = 226;
// bram[29152] = 215;
// bram[29153] = 201;
// bram[29154] = 187;
// bram[29155] = 171;
// bram[29156] = 154;
// bram[29157] = 137;
// bram[29158] = 119;
// bram[29159] = 102;
// bram[29160] = 85;
// bram[29161] = 69;
// bram[29162] = 54;
// bram[29163] = 41;
// bram[29164] = 29;
// bram[29165] = 19;
// bram[29166] = 10;
// bram[29167] = 5;
// bram[29168] = 1;
// bram[29169] = 0;
// bram[29170] = 1;
// bram[29171] = 4;
// bram[29172] = 10;
// bram[29173] = 18;
// bram[29174] = 28;
// bram[29175] = 39;
// bram[29176] = 53;
// bram[29177] = 68;
// bram[29178] = 84;
// bram[29179] = 100;
// bram[29180] = 118;
// bram[29181] = 135;
// bram[29182] = 152;
// bram[29183] = 169;
// bram[29184] = 185;
// bram[29185] = 200;
// bram[29186] = 213;
// bram[29187] = 225;
// bram[29188] = 235;
// bram[29189] = 243;
// bram[29190] = 249;
// bram[29191] = 252;
// bram[29192] = 253;
// bram[29193] = 252;
// bram[29194] = 249;
// bram[29195] = 243;
// bram[29196] = 235;
// bram[29197] = 225;
// bram[29198] = 213;
// bram[29199] = 199;
// bram[29200] = 184;
// bram[29201] = 168;
// bram[29202] = 151;
// bram[29203] = 134;
// bram[29204] = 117;
// bram[29205] = 100;
// bram[29206] = 83;
// bram[29207] = 67;
// bram[29208] = 52;
// bram[29209] = 39;
// bram[29210] = 27;
// bram[29211] = 17;
// bram[29212] = 9;
// bram[29213] = 4;
// bram[29214] = 0;
// bram[29215] = 0;
// bram[29216] = 1;
// bram[29217] = 5;
// bram[29218] = 11;
// bram[29219] = 19;
// bram[29220] = 29;
// bram[29221] = 41;
// bram[29222] = 55;
// bram[29223] = 70;
// bram[29224] = 86;
// bram[29225] = 103;
// bram[29226] = 120;
// bram[29227] = 138;
// bram[29228] = 155;
// bram[29229] = 171;
// bram[29230] = 187;
// bram[29231] = 202;
// bram[29232] = 215;
// bram[29233] = 227;
// bram[29234] = 236;
// bram[29235] = 244;
// bram[29236] = 250;
// bram[29237] = 253;
// bram[29238] = 253;
// bram[29239] = 252;
// bram[29240] = 248;
// bram[29241] = 242;
// bram[29242] = 233;
// bram[29243] = 223;
// bram[29244] = 211;
// bram[29245] = 197;
// bram[29246] = 182;
// bram[29247] = 166;
// bram[29248] = 149;
// bram[29249] = 131;
// bram[29250] = 114;
// bram[29251] = 97;
// bram[29252] = 80;
// bram[29253] = 65;
// bram[29254] = 50;
// bram[29255] = 37;
// bram[29256] = 25;
// bram[29257] = 16;
// bram[29258] = 8;
// bram[29259] = 3;
// bram[29260] = 0;
// bram[29261] = 0;
// bram[29262] = 1;
// bram[29263] = 6;
// bram[29264] = 12;
// bram[29265] = 20;
// bram[29266] = 31;
// bram[29267] = 43;
// bram[29268] = 57;
// bram[29269] = 72;
// bram[29270] = 89;
// bram[29271] = 106;
// bram[29272] = 123;
// bram[29273] = 140;
// bram[29274] = 157;
// bram[29275] = 174;
// bram[29276] = 190;
// bram[29277] = 204;
// bram[29278] = 217;
// bram[29279] = 228;
// bram[29280] = 238;
// bram[29281] = 245;
// bram[29282] = 250;
// bram[29283] = 253;
// bram[29284] = 253;
// bram[29285] = 251;
// bram[29286] = 247;
// bram[29287] = 240;
// bram[29288] = 232;
// bram[29289] = 221;
// bram[29290] = 209;
// bram[29291] = 195;
// bram[29292] = 179;
// bram[29293] = 163;
// bram[29294] = 146;
// bram[29295] = 129;
// bram[29296] = 111;
// bram[29297] = 94;
// bram[29298] = 78;
// bram[29299] = 62;
// bram[29300] = 48;
// bram[29301] = 35;
// bram[29302] = 24;
// bram[29303] = 15;
// bram[29304] = 7;
// bram[29305] = 3;
// bram[29306] = 0;
// bram[29307] = 0;
// bram[29308] = 2;
// bram[29309] = 6;
// bram[29310] = 13;
// bram[29311] = 22;
// bram[29312] = 33;
// bram[29313] = 45;
// bram[29314] = 60;
// bram[29315] = 75;
// bram[29316] = 91;
// bram[29317] = 108;
// bram[29318] = 126;
// bram[29319] = 143;
// bram[29320] = 160;
// bram[29321] = 176;
// bram[29322] = 192;
// bram[29323] = 206;
// bram[29324] = 219;
// bram[29325] = 230;
// bram[29326] = 239;
// bram[29327] = 246;
// bram[29328] = 251;
// bram[29329] = 253;
// bram[29330] = 253;
// bram[29331] = 251;
// bram[29332] = 246;
// bram[29333] = 239;
// bram[29334] = 230;
// bram[29335] = 219;
// bram[29336] = 207;
// bram[29337] = 192;
// bram[29338] = 177;
// bram[29339] = 160;
// bram[29340] = 143;
// bram[29341] = 126;
// bram[29342] = 109;
// bram[29343] = 92;
// bram[29344] = 75;
// bram[29345] = 60;
// bram[29346] = 46;
// bram[29347] = 33;
// bram[29348] = 22;
// bram[29349] = 13;
// bram[29350] = 7;
// bram[29351] = 2;
// bram[29352] = 0;
// bram[29353] = 0;
// bram[29354] = 2;
// bram[29355] = 7;
// bram[29356] = 14;
// bram[29357] = 24;
// bram[29358] = 35;
// bram[29359] = 48;
// bram[29360] = 62;
// bram[29361] = 77;
// bram[29362] = 94;
// bram[29363] = 111;
// bram[29364] = 128;
// bram[29365] = 146;
// bram[29366] = 163;
// bram[29367] = 179;
// bram[29368] = 194;
// bram[29369] = 208;
// bram[29370] = 221;
// bram[29371] = 232;
// bram[29372] = 240;
// bram[29373] = 247;
// bram[29374] = 251;
// bram[29375] = 253;
// bram[29376] = 253;
// bram[29377] = 250;
// bram[29378] = 245;
// bram[29379] = 238;
// bram[29380] = 229;
// bram[29381] = 217;
// bram[29382] = 204;
// bram[29383] = 190;
// bram[29384] = 174;
// bram[29385] = 158;
// bram[29386] = 141;
// bram[29387] = 123;
// bram[29388] = 106;
// bram[29389] = 89;
// bram[29390] = 73;
// bram[29391] = 58;
// bram[29392] = 44;
// bram[29393] = 31;
// bram[29394] = 21;
// bram[29395] = 12;
// bram[29396] = 6;
// bram[29397] = 1;
// bram[29398] = 0;
// bram[29399] = 0;
// bram[29400] = 3;
// bram[29401] = 8;
// bram[29402] = 16;
// bram[29403] = 25;
// bram[29404] = 37;
// bram[29405] = 50;
// bram[29406] = 64;
// bram[29407] = 80;
// bram[29408] = 96;
// bram[29409] = 114;
// bram[29410] = 131;
// bram[29411] = 148;
// bram[29412] = 165;
// bram[29413] = 181;
// bram[29414] = 196;
// bram[29415] = 210;
// bram[29416] = 223;
// bram[29417] = 233;
// bram[29418] = 241;
// bram[29419] = 248;
// bram[29420] = 252;
// bram[29421] = 253;
// bram[29422] = 253;
// bram[29423] = 250;
// bram[29424] = 244;
// bram[29425] = 237;
// bram[29426] = 227;
// bram[29427] = 215;
// bram[29428] = 202;
// bram[29429] = 188;
// bram[29430] = 172;
// bram[29431] = 155;
// bram[29432] = 138;
// bram[29433] = 121;
// bram[29434] = 103;
// bram[29435] = 87;
// bram[29436] = 70;
// bram[29437] = 55;
// bram[29438] = 42;
// bram[29439] = 30;
// bram[29440] = 19;
// bram[29441] = 11;
// bram[29442] = 5;
// bram[29443] = 1;
// bram[29444] = 0;
// bram[29445] = 0;
// bram[29446] = 4;
// bram[29447] = 9;
// bram[29448] = 17;
// bram[29449] = 27;
// bram[29450] = 38;
// bram[29451] = 52;
// bram[29452] = 67;
// bram[29453] = 82;
// bram[29454] = 99;
// bram[29455] = 116;
// bram[29456] = 134;
// bram[29457] = 151;
// bram[29458] = 168;
// bram[29459] = 184;
// bram[29460] = 199;
// bram[29461] = 212;
// bram[29462] = 224;
// bram[29463] = 234;
// bram[29464] = 243;
// bram[29465] = 249;
// bram[29466] = 252;
// bram[29467] = 253;
// bram[29468] = 252;
// bram[29469] = 249;
// bram[29470] = 243;
// bram[29471] = 235;
// bram[29472] = 225;
// bram[29473] = 214;
// bram[29474] = 200;
// bram[29475] = 185;
// bram[29476] = 169;
// bram[29477] = 153;
// bram[29478] = 135;
// bram[29479] = 118;
// bram[29480] = 101;
// bram[29481] = 84;
// bram[29482] = 68;
// bram[29483] = 53;
// bram[29484] = 40;
// bram[29485] = 28;
// bram[29486] = 18;
// bram[29487] = 10;
// bram[29488] = 4;
// bram[29489] = 1;
// bram[29490] = 0;
// bram[29491] = 1;
// bram[29492] = 4;
// bram[29493] = 10;
// bram[29494] = 18;
// bram[29495] = 28;
// bram[29496] = 40;
// bram[29497] = 54;
// bram[29498] = 69;
// bram[29499] = 85;
// bram[29500] = 102;
// bram[29501] = 119;
// bram[29502] = 136;
// bram[29503] = 154;
// bram[29504] = 170;
// bram[29505] = 186;
// bram[29506] = 201;
// bram[29507] = 214;
// bram[29508] = 226;
// bram[29509] = 236;
// bram[29510] = 244;
// bram[29511] = 249;
// bram[29512] = 253;
// bram[29513] = 253;
// bram[29514] = 252;
// bram[29515] = 248;
// bram[29516] = 242;
// bram[29517] = 234;
// bram[29518] = 224;
// bram[29519] = 212;
// bram[29520] = 198;
// bram[29521] = 183;
// bram[29522] = 167;
// bram[29523] = 150;
// bram[29524] = 133;
// bram[29525] = 115;
// bram[29526] = 98;
// bram[29527] = 81;
// bram[29528] = 66;
// bram[29529] = 51;
// bram[29530] = 38;
// bram[29531] = 26;
// bram[29532] = 16;
// bram[29533] = 9;
// bram[29534] = 3;
// bram[29535] = 0;
// bram[29536] = 0;
// bram[29537] = 1;
// bram[29538] = 5;
// bram[29539] = 11;
// bram[29540] = 20;
// bram[29541] = 30;
// bram[29542] = 42;
// bram[29543] = 56;
// bram[29544] = 71;
// bram[29545] = 87;
// bram[29546] = 104;
// bram[29547] = 122;
// bram[29548] = 139;
// bram[29549] = 156;
// bram[29550] = 173;
// bram[29551] = 189;
// bram[29552] = 203;
// bram[29553] = 216;
// bram[29554] = 228;
// bram[29555] = 237;
// bram[29556] = 245;
// bram[29557] = 250;
// bram[29558] = 253;
// bram[29559] = 253;
// bram[29560] = 252;
// bram[29561] = 247;
// bram[29562] = 241;
// bram[29563] = 232;
// bram[29564] = 222;
// bram[29565] = 210;
// bram[29566] = 196;
// bram[29567] = 180;
// bram[29568] = 164;
// bram[29569] = 147;
// bram[29570] = 130;
// bram[29571] = 113;
// bram[29572] = 95;
// bram[29573] = 79;
// bram[29574] = 63;
// bram[29575] = 49;
// bram[29576] = 36;
// bram[29577] = 25;
// bram[29578] = 15;
// bram[29579] = 8;
// bram[29580] = 3;
// bram[29581] = 0;
// bram[29582] = 0;
// bram[29583] = 2;
// bram[29584] = 6;
// bram[29585] = 13;
// bram[29586] = 21;
// bram[29587] = 32;
// bram[29588] = 44;
// bram[29589] = 58;
// bram[29590] = 74;
// bram[29591] = 90;
// bram[29592] = 107;
// bram[29593] = 124;
// bram[29594] = 142;
// bram[29595] = 159;
// bram[29596] = 175;
// bram[29597] = 191;
// bram[29598] = 205;
// bram[29599] = 218;
// bram[29600] = 229;
// bram[29601] = 238;
// bram[29602] = 246;
// bram[29603] = 251;
// bram[29604] = 253;
// bram[29605] = 253;
// bram[29606] = 251;
// bram[29607] = 247;
// bram[29608] = 240;
// bram[29609] = 231;
// bram[29610] = 220;
// bram[29611] = 207;
// bram[29612] = 193;
// bram[29613] = 178;
// bram[29614] = 162;
// bram[29615] = 145;
// bram[29616] = 127;
// bram[29617] = 110;
// bram[29618] = 93;
// bram[29619] = 76;
// bram[29620] = 61;
// bram[29621] = 47;
// bram[29622] = 34;
// bram[29623] = 23;
// bram[29624] = 14;
// bram[29625] = 7;
// bram[29626] = 2;
// bram[29627] = 0;
// bram[29628] = 0;
// bram[29629] = 2;
// bram[29630] = 7;
// bram[29631] = 14;
// bram[29632] = 23;
// bram[29633] = 34;
// bram[29634] = 47;
// bram[29635] = 61;
// bram[29636] = 76;
// bram[29637] = 93;
// bram[29638] = 110;
// bram[29639] = 127;
// bram[29640] = 144;
// bram[29641] = 161;
// bram[29642] = 178;
// bram[29643] = 193;
// bram[29644] = 207;
// bram[29645] = 220;
// bram[29646] = 231;
// bram[29647] = 240;
// bram[29648] = 247;
// bram[29649] = 251;
// bram[29650] = 253;
// bram[29651] = 253;
// bram[29652] = 251;
// bram[29653] = 246;
// bram[29654] = 239;
// bram[29655] = 229;
// bram[29656] = 218;
// bram[29657] = 205;
// bram[29658] = 191;
// bram[29659] = 176;
// bram[29660] = 159;
// bram[29661] = 142;
// bram[29662] = 125;
// bram[29663] = 107;
// bram[29664] = 90;
// bram[29665] = 74;
// bram[29666] = 59;
// bram[29667] = 45;
// bram[29668] = 32;
// bram[29669] = 21;
// bram[29670] = 13;
// bram[29671] = 6;
// bram[29672] = 2;
// bram[29673] = 0;
// bram[29674] = 0;
// bram[29675] = 3;
// bram[29676] = 8;
// bram[29677] = 15;
// bram[29678] = 24;
// bram[29679] = 36;
// bram[29680] = 49;
// bram[29681] = 63;
// bram[29682] = 79;
// bram[29683] = 95;
// bram[29684] = 112;
// bram[29685] = 130;
// bram[29686] = 147;
// bram[29687] = 164;
// bram[29688] = 180;
// bram[29689] = 195;
// bram[29690] = 209;
// bram[29691] = 222;
// bram[29692] = 232;
// bram[29693] = 241;
// bram[29694] = 247;
// bram[29695] = 252;
// bram[29696] = 253;
// bram[29697] = 253;
// bram[29698] = 250;
// bram[29699] = 245;
// bram[29700] = 237;
// bram[29701] = 228;
// bram[29702] = 216;
// bram[29703] = 203;
// bram[29704] = 189;
// bram[29705] = 173;
// bram[29706] = 156;
// bram[29707] = 139;
// bram[29708] = 122;
// bram[29709] = 105;
// bram[29710] = 88;
// bram[29711] = 72;
// bram[29712] = 56;
// bram[29713] = 43;
// bram[29714] = 30;
// bram[29715] = 20;
// bram[29716] = 12;
// bram[29717] = 5;
// bram[29718] = 1;
// bram[29719] = 0;
// bram[29720] = 0;
// bram[29721] = 3;
// bram[29722] = 9;
// bram[29723] = 16;
// bram[29724] = 26;
// bram[29725] = 38;
// bram[29726] = 51;
// bram[29727] = 65;
// bram[29728] = 81;
// bram[29729] = 98;
// bram[29730] = 115;
// bram[29731] = 132;
// bram[29732] = 150;
// bram[29733] = 167;
// bram[29734] = 183;
// bram[29735] = 198;
// bram[29736] = 211;
// bram[29737] = 223;
// bram[29738] = 234;
// bram[29739] = 242;
// bram[29740] = 248;
// bram[29741] = 252;
// bram[29742] = 253;
// bram[29743] = 253;
// bram[29744] = 249;
// bram[29745] = 244;
// bram[29746] = 236;
// bram[29747] = 226;
// bram[29748] = 214;
// bram[29749] = 201;
// bram[29750] = 186;
// bram[29751] = 171;
// bram[29752] = 154;
// bram[29753] = 137;
// bram[29754] = 119;
// bram[29755] = 102;
// bram[29756] = 85;
// bram[29757] = 69;
// bram[29758] = 54;
// bram[29759] = 41;
// bram[29760] = 29;
// bram[29761] = 19;
// bram[29762] = 10;
// bram[29763] = 4;
// bram[29764] = 1;
// bram[29765] = 0;
// bram[29766] = 1;
// bram[29767] = 4;
// bram[29768] = 10;
// bram[29769] = 18;
// bram[29770] = 28;
// bram[29771] = 40;
// bram[29772] = 53;
// bram[29773] = 68;
// bram[29774] = 84;
// bram[29775] = 101;
// bram[29776] = 118;
// bram[29777] = 135;
// bram[29778] = 152;
// bram[29779] = 169;
// bram[29780] = 185;
// bram[29781] = 200;
// bram[29782] = 213;
// bram[29783] = 225;
// bram[29784] = 235;
// bram[29785] = 243;
// bram[29786] = 249;
// bram[29787] = 252;
// bram[29788] = 253;
// bram[29789] = 252;
// bram[29790] = 249;
// bram[29791] = 243;
// bram[29792] = 235;
// bram[29793] = 224;
// bram[29794] = 212;
// bram[29795] = 199;
// bram[29796] = 184;
// bram[29797] = 168;
// bram[29798] = 151;
// bram[29799] = 134;
// bram[29800] = 117;
// bram[29801] = 99;
// bram[29802] = 83;
// bram[29803] = 67;
// bram[29804] = 52;
// bram[29805] = 39;
// bram[29806] = 27;
// bram[29807] = 17;
// bram[29808] = 9;
// bram[29809] = 4;
// bram[29810] = 0;
// bram[29811] = 0;
// bram[29812] = 1;
// bram[29813] = 5;
// bram[29814] = 11;
// bram[29815] = 19;
// bram[29816] = 29;
// bram[29817] = 42;
// bram[29818] = 55;
// bram[29819] = 70;
// bram[29820] = 86;
// bram[29821] = 103;
// bram[29822] = 120;
// bram[29823] = 138;
// bram[29824] = 155;
// bram[29825] = 172;
// bram[29826] = 187;
// bram[29827] = 202;
// bram[29828] = 215;
// bram[29829] = 227;
// bram[29830] = 237;
// bram[29831] = 244;
// bram[29832] = 250;
// bram[29833] = 253;
// bram[29834] = 253;
// bram[29835] = 252;
// bram[29836] = 248;
// bram[29837] = 242;
// bram[29838] = 233;
// bram[29839] = 223;
// bram[29840] = 210;
// bram[29841] = 197;
// bram[29842] = 182;
// bram[29843] = 165;
// bram[29844] = 149;
// bram[29845] = 131;
// bram[29846] = 114;
// bram[29847] = 97;
// bram[29848] = 80;
// bram[29849] = 64;
// bram[29850] = 50;
// bram[29851] = 37;
// bram[29852] = 25;
// bram[29853] = 16;
// bram[29854] = 8;
// bram[29855] = 3;
// bram[29856] = 0;
// bram[29857] = 0;
// bram[29858] = 1;
// bram[29859] = 6;
// bram[29860] = 12;
// bram[29861] = 21;
// bram[29862] = 31;
// bram[29863] = 44;
// bram[29864] = 57;
// bram[29865] = 73;
// bram[29866] = 89;
// bram[29867] = 106;
// bram[29868] = 123;
// bram[29869] = 140;
// bram[29870] = 158;
// bram[29871] = 174;
// bram[29872] = 190;
// bram[29873] = 204;
// bram[29874] = 217;
// bram[29875] = 229;
// bram[29876] = 238;
// bram[29877] = 245;
// bram[29878] = 250;
// bram[29879] = 253;
// bram[29880] = 253;
// bram[29881] = 251;
// bram[29882] = 247;
// bram[29883] = 240;
// bram[29884] = 232;
// bram[29885] = 221;
// bram[29886] = 208;
// bram[29887] = 194;
// bram[29888] = 179;
// bram[29889] = 163;
// bram[29890] = 146;
// bram[29891] = 129;
// bram[29892] = 111;
// bram[29893] = 94;
// bram[29894] = 78;
// bram[29895] = 62;
// bram[29896] = 48;
// bram[29897] = 35;
// bram[29898] = 24;
// bram[29899] = 14;
// bram[29900] = 7;
// bram[29901] = 2;
// bram[29902] = 0;
// bram[29903] = 0;
// bram[29904] = 2;
// bram[29905] = 6;
// bram[29906] = 13;
// bram[29907] = 22;
// bram[29908] = 33;
// bram[29909] = 46;
// bram[29910] = 60;
// bram[29911] = 75;
// bram[29912] = 91;
// bram[29913] = 108;
// bram[29914] = 126;
// bram[29915] = 143;
// bram[29916] = 160;
// bram[29917] = 177;
// bram[29918] = 192;
// bram[29919] = 206;
// bram[29920] = 219;
// bram[29921] = 230;
// bram[29922] = 239;
// bram[29923] = 246;
// bram[29924] = 251;
// bram[29925] = 253;
// bram[29926] = 253;
// bram[29927] = 251;
// bram[29928] = 246;
// bram[29929] = 239;
// bram[29930] = 230;
// bram[29931] = 219;
// bram[29932] = 206;
// bram[29933] = 192;
// bram[29934] = 177;
// bram[29935] = 160;
// bram[29936] = 143;
// bram[29937] = 126;
// bram[29938] = 109;
// bram[29939] = 91;
// bram[29940] = 75;
// bram[29941] = 60;
// bram[29942] = 46;
// bram[29943] = 33;
// bram[29944] = 22;
// bram[29945] = 13;
// bram[29946] = 6;
// bram[29947] = 2;
// bram[29948] = 0;
// bram[29949] = 0;
// bram[29950] = 2;
// bram[29951] = 7;
// bram[29952] = 14;
// bram[29953] = 24;
// bram[29954] = 35;
// bram[29955] = 48;
// bram[29956] = 62;
// bram[29957] = 78;
// bram[29958] = 94;
// bram[29959] = 111;
// bram[29960] = 128;
// bram[29961] = 146;
// bram[29962] = 163;
// bram[29963] = 179;
// bram[29964] = 194;
// bram[29965] = 208;
// bram[29966] = 221;
// bram[29967] = 232;
// bram[29968] = 240;
// bram[29969] = 247;
// bram[29970] = 251;
// bram[29971] = 253;
// bram[29972] = 253;
// bram[29973] = 250;
// bram[29974] = 245;
// bram[29975] = 238;
// bram[29976] = 229;
// bram[29977] = 217;
// bram[29978] = 204;
// bram[29979] = 190;
// bram[29980] = 174;
// bram[29981] = 158;
// bram[29982] = 141;
// bram[29983] = 123;
// bram[29984] = 106;
// bram[29985] = 89;
// bram[29986] = 73;
// bram[29987] = 57;
// bram[29988] = 44;
// bram[29989] = 31;
// bram[29990] = 21;
// bram[29991] = 12;
// bram[29992] = 6;
// bram[29993] = 1;
// bram[29994] = 0;
// bram[29995] = 0;
// bram[29996] = 3;
// bram[29997] = 8;
// bram[29998] = 16;
// bram[29999] = 25;
// bram[30000] = 37;
// bram[30001] = 50;
// bram[30002] = 64;
// bram[30003] = 80;
// bram[30004] = 97;
// bram[30005] = 114;
// bram[30006] = 131;
// bram[30007] = 148;
// bram[30008] = 165;
// bram[30009] = 182;
// bram[30010] = 197;
// bram[30011] = 210;
// bram[30012] = 223;
// bram[30013] = 233;
// bram[30014] = 242;
// bram[30015] = 248;
// bram[30016] = 252;
// bram[30017] = 253;
// bram[30018] = 253;
// bram[30019] = 250;
// bram[30020] = 244;
// bram[30021] = 237;
// bram[30022] = 227;
// bram[30023] = 215;
// bram[30024] = 202;
// bram[30025] = 187;
// bram[30026] = 172;
// bram[30027] = 155;
// bram[30028] = 138;
// bram[30029] = 120;
// bram[30030] = 103;
// bram[30031] = 86;
// bram[30032] = 70;
// bram[30033] = 55;
// bram[30034] = 42;
// bram[30035] = 29;
// bram[30036] = 19;
// bram[30037] = 11;
// bram[30038] = 5;
// bram[30039] = 1;
// bram[30040] = 0;
// bram[30041] = 0;
// bram[30042] = 4;
// bram[30043] = 9;
// bram[30044] = 17;
// bram[30045] = 27;
// bram[30046] = 39;
// bram[30047] = 52;
// bram[30048] = 67;
// bram[30049] = 83;
// bram[30050] = 99;
// bram[30051] = 116;
// bram[30052] = 134;
// bram[30053] = 151;
// bram[30054] = 168;
// bram[30055] = 184;
// bram[30056] = 199;
// bram[30057] = 212;
// bram[30058] = 224;
// bram[30059] = 235;
// bram[30060] = 243;
// bram[30061] = 249;
// bram[30062] = 252;
// bram[30063] = 253;
// bram[30064] = 252;
// bram[30065] = 249;
// bram[30066] = 243;
// bram[30067] = 235;
// bram[30068] = 225;
// bram[30069] = 213;
// bram[30070] = 200;
// bram[30071] = 185;
// bram[30072] = 169;
// bram[30073] = 152;
// bram[30074] = 135;
// bram[30075] = 118;
// bram[30076] = 101;
// bram[30077] = 84;
// bram[30078] = 68;
// bram[30079] = 53;
// bram[30080] = 40;
// bram[30081] = 28;
// bram[30082] = 18;
// bram[30083] = 10;
// bram[30084] = 4;
// bram[30085] = 1;
// bram[30086] = 0;
// bram[30087] = 1;
// bram[30088] = 4;
// bram[30089] = 10;
// bram[30090] = 18;
// bram[30091] = 29;
// bram[30092] = 41;
// bram[30093] = 54;
// bram[30094] = 69;
// bram[30095] = 85;
// bram[30096] = 102;
// bram[30097] = 119;
// bram[30098] = 137;
// bram[30099] = 154;
// bram[30100] = 170;
// bram[30101] = 186;
// bram[30102] = 201;
// bram[30103] = 214;
// bram[30104] = 226;
// bram[30105] = 236;
// bram[30106] = 244;
// bram[30107] = 249;
// bram[30108] = 253;
// bram[30109] = 253;
// bram[30110] = 252;
// bram[30111] = 248;
// bram[30112] = 242;
// bram[30113] = 234;
// bram[30114] = 224;
// bram[30115] = 211;
// bram[30116] = 198;
// bram[30117] = 183;
// bram[30118] = 167;
// bram[30119] = 150;
// bram[30120] = 132;
// bram[30121] = 115;
// bram[30122] = 98;
// bram[30123] = 81;
// bram[30124] = 65;
// bram[30125] = 51;
// bram[30126] = 38;
// bram[30127] = 26;
// bram[30128] = 16;
// bram[30129] = 9;
// bram[30130] = 3;
// bram[30131] = 0;
// bram[30132] = 0;
// bram[30133] = 1;
// bram[30134] = 5;
// bram[30135] = 11;
// bram[30136] = 20;
// bram[30137] = 30;
// bram[30138] = 43;
// bram[30139] = 56;
// bram[30140] = 72;
// bram[30141] = 88;
// bram[30142] = 105;
// bram[30143] = 122;
// bram[30144] = 139;
// bram[30145] = 156;
// bram[30146] = 173;
// bram[30147] = 189;
// bram[30148] = 203;
// bram[30149] = 216;
// bram[30150] = 228;
// bram[30151] = 237;
// bram[30152] = 245;
// bram[30153] = 250;
// bram[30154] = 253;
// bram[30155] = 253;
// bram[30156] = 252;
// bram[30157] = 247;
// bram[30158] = 241;
// bram[30159] = 232;
// bram[30160] = 222;
// bram[30161] = 209;
// bram[30162] = 195;
// bram[30163] = 180;
// bram[30164] = 164;
// bram[30165] = 147;
// bram[30166] = 130;
// bram[30167] = 112;
// bram[30168] = 95;
// bram[30169] = 79;
// bram[30170] = 63;
// bram[30171] = 49;
// bram[30172] = 36;
// bram[30173] = 24;
// bram[30174] = 15;
// bram[30175] = 8;
// bram[30176] = 3;
// bram[30177] = 0;
// bram[30178] = 0;
// bram[30179] = 2;
// bram[30180] = 6;
// bram[30181] = 13;
// bram[30182] = 21;
// bram[30183] = 32;
// bram[30184] = 45;
// bram[30185] = 59;
// bram[30186] = 74;
// bram[30187] = 90;
// bram[30188] = 107;
// bram[30189] = 125;
// bram[30190] = 142;
// bram[30191] = 159;
// bram[30192] = 175;
// bram[30193] = 191;
// bram[30194] = 205;
// bram[30195] = 218;
// bram[30196] = 229;
// bram[30197] = 239;
// bram[30198] = 246;
// bram[30199] = 251;
// bram[30200] = 253;
// bram[30201] = 253;
// bram[30202] = 251;
// bram[30203] = 247;
// bram[30204] = 240;
// bram[30205] = 231;
// bram[30206] = 220;
// bram[30207] = 207;
// bram[30208] = 193;
// bram[30209] = 178;
// bram[30210] = 161;
// bram[30211] = 144;
// bram[30212] = 127;
// bram[30213] = 110;
// bram[30214] = 93;
// bram[30215] = 76;
// bram[30216] = 61;
// bram[30217] = 47;
// bram[30218] = 34;
// bram[30219] = 23;
// bram[30220] = 14;
// bram[30221] = 7;
// bram[30222] = 2;
// bram[30223] = 0;
// bram[30224] = 0;
// bram[30225] = 2;
// bram[30226] = 7;
// bram[30227] = 14;
// bram[30228] = 23;
// bram[30229] = 34;
// bram[30230] = 47;
// bram[30231] = 61;
// bram[30232] = 76;
// bram[30233] = 93;
// bram[30234] = 110;
// bram[30235] = 127;
// bram[30236] = 145;
// bram[30237] = 162;
// bram[30238] = 178;
// bram[30239] = 193;
// bram[30240] = 207;
// bram[30241] = 220;
// bram[30242] = 231;
// bram[30243] = 240;
// bram[30244] = 247;
// bram[30245] = 251;
// bram[30246] = 253;
// bram[30247] = 253;
// bram[30248] = 251;
// bram[30249] = 246;
// bram[30250] = 239;
// bram[30251] = 229;
// bram[30252] = 218;
// bram[30253] = 205;
// bram[30254] = 191;
// bram[30255] = 175;
// bram[30256] = 159;
// bram[30257] = 142;
// bram[30258] = 124;
// bram[30259] = 107;
// bram[30260] = 90;
// bram[30261] = 74;
// bram[30262] = 59;
// bram[30263] = 45;
// bram[30264] = 32;
// bram[30265] = 21;
// bram[30266] = 13;
// bram[30267] = 6;
// bram[30268] = 2;
// bram[30269] = 0;
// bram[30270] = 0;
// bram[30271] = 3;
// bram[30272] = 8;
// bram[30273] = 15;
// bram[30274] = 25;
// bram[30275] = 36;
// bram[30276] = 49;
// bram[30277] = 63;
// bram[30278] = 79;
// bram[30279] = 95;
// bram[30280] = 113;
// bram[30281] = 130;
// bram[30282] = 147;
// bram[30283] = 164;
// bram[30284] = 180;
// bram[30285] = 196;
// bram[30286] = 210;
// bram[30287] = 222;
// bram[30288] = 232;
// bram[30289] = 241;
// bram[30290] = 247;
// bram[30291] = 252;
// bram[30292] = 253;
// bram[30293] = 253;
// bram[30294] = 250;
// bram[30295] = 245;
// bram[30296] = 237;
// bram[30297] = 228;
// bram[30298] = 216;
// bram[30299] = 203;
// bram[30300] = 189;
// bram[30301] = 173;
// bram[30302] = 156;
// bram[30303] = 139;
// bram[30304] = 122;
// bram[30305] = 104;
// bram[30306] = 88;
// bram[30307] = 71;
// bram[30308] = 56;
// bram[30309] = 42;
// bram[30310] = 30;
// bram[30311] = 20;
// bram[30312] = 11;
// bram[30313] = 5;
// bram[30314] = 1;
// bram[30315] = 0;
// bram[30316] = 0;
// bram[30317] = 3;
// bram[30318] = 9;
// bram[30319] = 16;
// bram[30320] = 26;
// bram[30321] = 38;
// bram[30322] = 51;
// bram[30323] = 66;
// bram[30324] = 81;
// bram[30325] = 98;
// bram[30326] = 115;
// bram[30327] = 133;
// bram[30328] = 150;
// bram[30329] = 167;
// bram[30330] = 183;
// bram[30331] = 198;
// bram[30332] = 212;
// bram[30333] = 224;
// bram[30334] = 234;
// bram[30335] = 242;
// bram[30336] = 248;
// bram[30337] = 252;
// bram[30338] = 253;
// bram[30339] = 253;
// bram[30340] = 249;
// bram[30341] = 244;
// bram[30342] = 236;
// bram[30343] = 226;
// bram[30344] = 214;
// bram[30345] = 201;
// bram[30346] = 186;
// bram[30347] = 170;
// bram[30348] = 154;
// bram[30349] = 136;
// bram[30350] = 119;
// bram[30351] = 102;
// bram[30352] = 85;
// bram[30353] = 69;
// bram[30354] = 54;
// bram[30355] = 40;
// bram[30356] = 29;
// bram[30357] = 18;
// bram[30358] = 10;
// bram[30359] = 4;
// bram[30360] = 1;
// bram[30361] = 0;
// bram[30362] = 1;
// bram[30363] = 4;
// bram[30364] = 10;
// bram[30365] = 18;
// bram[30366] = 28;
// bram[30367] = 40;
// bram[30368] = 53;
// bram[30369] = 68;
// bram[30370] = 84;
// bram[30371] = 101;
// bram[30372] = 118;
// bram[30373] = 135;
// bram[30374] = 153;
// bram[30375] = 169;
// bram[30376] = 185;
// bram[30377] = 200;
// bram[30378] = 214;
// bram[30379] = 225;
// bram[30380] = 235;
// bram[30381] = 243;
// bram[30382] = 249;
// bram[30383] = 252;
// bram[30384] = 253;
// bram[30385] = 252;
// bram[30386] = 249;
// bram[30387] = 243;
// bram[30388] = 234;
// bram[30389] = 224;
// bram[30390] = 212;
// bram[30391] = 199;
// bram[30392] = 184;
// bram[30393] = 168;
// bram[30394] = 151;
// bram[30395] = 134;
// bram[30396] = 116;
// bram[30397] = 99;
// bram[30398] = 82;
// bram[30399] = 67;
// bram[30400] = 52;
// bram[30401] = 39;
// bram[30402] = 27;
// bram[30403] = 17;
// bram[30404] = 9;
// bram[30405] = 4;
// bram[30406] = 0;
// bram[30407] = 0;
// bram[30408] = 1;
// bram[30409] = 5;
// bram[30410] = 11;
// bram[30411] = 19;
// bram[30412] = 30;
// bram[30413] = 42;
// bram[30414] = 55;
// bram[30415] = 70;
// bram[30416] = 86;
// bram[30417] = 103;
// bram[30418] = 121;
// bram[30419] = 138;
// bram[30420] = 155;
// bram[30421] = 172;
// bram[30422] = 188;
// bram[30423] = 202;
// bram[30424] = 215;
// bram[30425] = 227;
// bram[30426] = 237;
// bram[30427] = 244;
// bram[30428] = 250;
// bram[30429] = 253;
// bram[30430] = 253;
// bram[30431] = 252;
// bram[30432] = 248;
// bram[30433] = 241;
// bram[30434] = 233;
// bram[30435] = 223;
// bram[30436] = 210;
// bram[30437] = 197;
// bram[30438] = 181;
// bram[30439] = 165;
// bram[30440] = 148;
// bram[30441] = 131;
// bram[30442] = 114;
// bram[30443] = 97;
// bram[30444] = 80;
// bram[30445] = 64;
// bram[30446] = 50;
// bram[30447] = 37;
// bram[30448] = 25;
// bram[30449] = 16;
// bram[30450] = 8;
// bram[30451] = 3;
// bram[30452] = 0;
// bram[30453] = 0;
// bram[30454] = 1;
// bram[30455] = 6;
// bram[30456] = 12;
// bram[30457] = 21;
// bram[30458] = 31;
// bram[30459] = 44;
// bram[30460] = 58;
// bram[30461] = 73;
// bram[30462] = 89;
// bram[30463] = 106;
// bram[30464] = 123;
// bram[30465] = 141;
// bram[30466] = 158;
// bram[30467] = 174;
// bram[30468] = 190;
// bram[30469] = 204;
// bram[30470] = 217;
// bram[30471] = 229;
// bram[30472] = 238;
// bram[30473] = 245;
// bram[30474] = 250;
// bram[30475] = 253;
// bram[30476] = 253;
// bram[30477] = 251;
// bram[30478] = 247;
// bram[30479] = 240;
// bram[30480] = 232;
// bram[30481] = 221;
// bram[30482] = 208;
// bram[30483] = 194;
// bram[30484] = 179;
// bram[30485] = 163;
// bram[30486] = 146;
// bram[30487] = 128;
// bram[30488] = 111;
// bram[30489] = 94;
// bram[30490] = 77;
// bram[30491] = 62;
// bram[30492] = 48;
// bram[30493] = 35;
// bram[30494] = 24;
// bram[30495] = 14;
// bram[30496] = 7;
// bram[30497] = 2;
// bram[30498] = 0;
// bram[30499] = 0;
// bram[30500] = 2;
// bram[30501] = 6;
// bram[30502] = 13;
// bram[30503] = 22;
// bram[30504] = 33;
// bram[30505] = 46;
// bram[30506] = 60;
// bram[30507] = 75;
// bram[30508] = 92;
// bram[30509] = 109;
// bram[30510] = 126;
// bram[30511] = 143;
// bram[30512] = 160;
// bram[30513] = 177;
// bram[30514] = 192;
// bram[30515] = 206;
// bram[30516] = 219;
// bram[30517] = 230;
// bram[30518] = 239;
// bram[30519] = 246;
// bram[30520] = 251;
// bram[30521] = 253;
// bram[30522] = 253;
// bram[30523] = 251;
// bram[30524] = 246;
// bram[30525] = 239;
// bram[30526] = 230;
// bram[30527] = 219;
// bram[30528] = 206;
// bram[30529] = 192;
// bram[30530] = 176;
// bram[30531] = 160;
// bram[30532] = 143;
// bram[30533] = 126;
// bram[30534] = 108;
// bram[30535] = 91;
// bram[30536] = 75;
// bram[30537] = 60;
// bram[30538] = 45;
// bram[30539] = 33;
// bram[30540] = 22;
// bram[30541] = 13;
// bram[30542] = 6;
// bram[30543] = 2;
// bram[30544] = 0;
// bram[30545] = 0;
// bram[30546] = 2;
// bram[30547] = 7;
// bram[30548] = 15;
// bram[30549] = 24;
// bram[30550] = 35;
// bram[30551] = 48;
// bram[30552] = 62;
// bram[30553] = 78;
// bram[30554] = 94;
// bram[30555] = 111;
// bram[30556] = 129;
// bram[30557] = 146;
// bram[30558] = 163;
// bram[30559] = 179;
// bram[30560] = 195;
// bram[30561] = 209;
// bram[30562] = 221;
// bram[30563] = 232;
// bram[30564] = 240;
// bram[30565] = 247;
// bram[30566] = 251;
// bram[30567] = 253;
// bram[30568] = 253;
// bram[30569] = 250;
// bram[30570] = 245;
// bram[30571] = 238;
// bram[30572] = 228;
// bram[30573] = 217;
// bram[30574] = 204;
// bram[30575] = 190;
// bram[30576] = 174;
// bram[30577] = 157;
// bram[30578] = 140;
// bram[30579] = 123;
// bram[30580] = 106;
// bram[30581] = 89;
// bram[30582] = 73;
// bram[30583] = 57;
// bram[30584] = 43;
// bram[30585] = 31;
// bram[30586] = 21;
// bram[30587] = 12;
// bram[30588] = 6;
// bram[30589] = 1;
// bram[30590] = 0;
// bram[30591] = 0;
// bram[30592] = 3;
// bram[30593] = 8;
// bram[30594] = 16;
// bram[30595] = 25;
// bram[30596] = 37;
// bram[30597] = 50;
// bram[30598] = 65;
// bram[30599] = 80;
// bram[30600] = 97;
// bram[30601] = 114;
// bram[30602] = 131;
// bram[30603] = 149;
// bram[30604] = 166;
// bram[30605] = 182;
// bram[30606] = 197;
// bram[30607] = 211;
// bram[30608] = 223;
// bram[30609] = 233;
// bram[30610] = 242;
// bram[30611] = 248;
// bram[30612] = 252;
// bram[30613] = 253;
// bram[30614] = 253;
// bram[30615] = 250;
// bram[30616] = 244;
// bram[30617] = 236;
// bram[30618] = 227;
// bram[30619] = 215;
// bram[30620] = 202;
// bram[30621] = 187;
// bram[30622] = 171;
// bram[30623] = 155;
// bram[30624] = 138;
// bram[30625] = 120;
// bram[30626] = 103;
// bram[30627] = 86;
// bram[30628] = 70;
// bram[30629] = 55;
// bram[30630] = 41;
// bram[30631] = 29;
// bram[30632] = 19;
// bram[30633] = 11;
// bram[30634] = 5;
// bram[30635] = 1;
// bram[30636] = 0;
// bram[30637] = 0;
// bram[30638] = 4;
// bram[30639] = 9;
// bram[30640] = 17;
// bram[30641] = 27;
// bram[30642] = 39;
// bram[30643] = 52;
// bram[30644] = 67;
// bram[30645] = 83;
// bram[30646] = 99;
// bram[30647] = 117;
// bram[30648] = 134;
// bram[30649] = 151;
// bram[30650] = 168;
// bram[30651] = 184;
// bram[30652] = 199;
// bram[30653] = 213;
// bram[30654] = 225;
// bram[30655] = 235;
// bram[30656] = 243;
// bram[30657] = 249;
// bram[30658] = 252;
// bram[30659] = 253;
// bram[30660] = 252;
// bram[30661] = 249;
// bram[30662] = 243;
// bram[30663] = 235;
// bram[30664] = 225;
// bram[30665] = 213;
// bram[30666] = 200;
// bram[30667] = 185;
// bram[30668] = 169;
// bram[30669] = 152;
// bram[30670] = 135;
// bram[30671] = 118;
// bram[30672] = 100;
// bram[30673] = 84;
// bram[30674] = 68;
// bram[30675] = 53;
// bram[30676] = 39;
// bram[30677] = 28;
// bram[30678] = 18;
// bram[30679] = 10;
// bram[30680] = 4;
// bram[30681] = 1;
// bram[30682] = 0;
// bram[30683] = 1;
// bram[30684] = 4;
// bram[30685] = 10;
// bram[30686] = 19;
// bram[30687] = 29;
// bram[30688] = 41;
// bram[30689] = 54;
// bram[30690] = 69;
// bram[30691] = 85;
// bram[30692] = 102;
// bram[30693] = 119;
// bram[30694] = 137;
// bram[30695] = 154;
// bram[30696] = 171;
// bram[30697] = 186;
// bram[30698] = 201;
// bram[30699] = 215;
// bram[30700] = 226;
// bram[30701] = 236;
// bram[30702] = 244;
// bram[30703] = 249;
// bram[30704] = 253;
// bram[30705] = 253;
// bram[30706] = 252;
// bram[30707] = 248;
// bram[30708] = 242;
// bram[30709] = 234;
// bram[30710] = 223;
// bram[30711] = 211;
// bram[30712] = 198;
// bram[30713] = 183;
// bram[30714] = 166;
// bram[30715] = 150;
// bram[30716] = 132;
// bram[30717] = 115;
// bram[30718] = 98;
// bram[30719] = 81;
// bram[30720] = 65;
// bram[30721] = 51;
// bram[30722] = 37;
// bram[30723] = 26;
// bram[30724] = 16;
// bram[30725] = 9;
// bram[30726] = 3;
// bram[30727] = 0;
// bram[30728] = 0;
// bram[30729] = 1;
// bram[30730] = 5;
// bram[30731] = 12;
// bram[30732] = 20;
// bram[30733] = 30;
// bram[30734] = 43;
// bram[30735] = 57;
// bram[30736] = 72;
// bram[30737] = 88;
// bram[30738] = 105;
// bram[30739] = 122;
// bram[30740] = 139;
// bram[30741] = 157;
// bram[30742] = 173;
// bram[30743] = 189;
// bram[30744] = 203;
// bram[30745] = 216;
// bram[30746] = 228;
// bram[30747] = 237;
// bram[30748] = 245;
// bram[30749] = 250;
// bram[30750] = 253;
// bram[30751] = 253;
// bram[30752] = 252;
// bram[30753] = 247;
// bram[30754] = 241;
// bram[30755] = 232;
// bram[30756] = 222;
// bram[30757] = 209;
// bram[30758] = 195;
// bram[30759] = 180;
// bram[30760] = 164;
// bram[30761] = 147;
// bram[30762] = 130;
// bram[30763] = 112;
// bram[30764] = 95;
// bram[30765] = 79;
// bram[30766] = 63;
// bram[30767] = 49;
// bram[30768] = 36;
// bram[30769] = 24;
// bram[30770] = 15;
// bram[30771] = 8;
// bram[30772] = 3;
// bram[30773] = 0;
// bram[30774] = 0;
// bram[30775] = 2;
// bram[30776] = 6;
// bram[30777] = 13;
// bram[30778] = 22;
// bram[30779] = 32;
// bram[30780] = 45;
// bram[30781] = 59;
// bram[30782] = 74;
// bram[30783] = 90;
// bram[30784] = 107;
// bram[30785] = 125;
// bram[30786] = 142;
// bram[30787] = 159;
// bram[30788] = 176;
// bram[30789] = 191;
// bram[30790] = 206;
// bram[30791] = 218;
// bram[30792] = 229;
// bram[30793] = 239;
// bram[30794] = 246;
// bram[30795] = 251;
// bram[30796] = 253;
// bram[30797] = 253;
// bram[30798] = 251;
// bram[30799] = 246;
// bram[30800] = 240;
// bram[30801] = 231;
// bram[30802] = 220;
// bram[30803] = 207;
// bram[30804] = 193;
// bram[30805] = 178;
// bram[30806] = 161;
// bram[30807] = 144;
// bram[30808] = 127;
// bram[30809] = 110;
// bram[30810] = 93;
// bram[30811] = 76;
// bram[30812] = 61;
// bram[30813] = 46;
// bram[30814] = 34;
// bram[30815] = 23;
// bram[30816] = 14;
// bram[30817] = 7;
// bram[30818] = 2;
// bram[30819] = 0;
// bram[30820] = 0;
// bram[30821] = 2;
// bram[30822] = 7;
// bram[30823] = 14;
// bram[30824] = 23;
// bram[30825] = 34;
// bram[30826] = 47;
// bram[30827] = 61;
// bram[30828] = 77;
// bram[30829] = 93;
// bram[30830] = 110;
// bram[30831] = 127;
// bram[30832] = 145;
// bram[30833] = 162;
// bram[30834] = 178;
// bram[30835] = 193;
// bram[30836] = 208;
// bram[30837] = 220;
// bram[30838] = 231;
// bram[30839] = 240;
// bram[30840] = 247;
// bram[30841] = 251;
// bram[30842] = 253;
// bram[30843] = 253;
// bram[30844] = 250;
// bram[30845] = 246;
// bram[30846] = 238;
// bram[30847] = 229;
// bram[30848] = 218;
// bram[30849] = 205;
// bram[30850] = 191;
// bram[30851] = 175;
// bram[30852] = 159;
// bram[30853] = 142;
// bram[30854] = 124;
// bram[30855] = 107;
// bram[30856] = 90;
// bram[30857] = 74;
// bram[30858] = 58;
// bram[30859] = 44;
// bram[30860] = 32;
// bram[30861] = 21;
// bram[30862] = 12;
// bram[30863] = 6;
// bram[30864] = 2;
// bram[30865] = 0;
// bram[30866] = 0;
// bram[30867] = 3;
// bram[30868] = 8;
// bram[30869] = 15;
// bram[30870] = 25;
// bram[30871] = 36;
// bram[30872] = 49;
// bram[30873] = 63;
// bram[30874] = 79;
// bram[30875] = 96;
// bram[30876] = 113;
// bram[30877] = 130;
// bram[30878] = 147;
// bram[30879] = 164;
// bram[30880] = 181;
// bram[30881] = 196;
// bram[30882] = 210;
// bram[30883] = 222;
// bram[30884] = 233;
// bram[30885] = 241;
// bram[30886] = 247;
// bram[30887] = 252;
// bram[30888] = 253;
// bram[30889] = 253;
// bram[30890] = 250;
// bram[30891] = 245;
// bram[30892] = 237;
// bram[30893] = 228;
// bram[30894] = 216;
// bram[30895] = 203;
// bram[30896] = 188;
// bram[30897] = 173;
// bram[30898] = 156;
// bram[30899] = 139;
// bram[30900] = 122;
// bram[30901] = 104;
// bram[30902] = 87;
// bram[30903] = 71;
// bram[30904] = 56;
// bram[30905] = 42;
// bram[30906] = 30;
// bram[30907] = 20;
// bram[30908] = 11;
// bram[30909] = 5;
// bram[30910] = 1;
// bram[30911] = 0;
// bram[30912] = 0;
// bram[30913] = 3;
// bram[30914] = 9;
// bram[30915] = 17;
// bram[30916] = 26;
// bram[30917] = 38;
// bram[30918] = 51;
// bram[30919] = 66;
// bram[30920] = 82;
// bram[30921] = 98;
// bram[30922] = 115;
// bram[30923] = 133;
// bram[30924] = 150;
// bram[30925] = 167;
// bram[30926] = 183;
// bram[30927] = 198;
// bram[30928] = 212;
// bram[30929] = 224;
// bram[30930] = 234;
// bram[30931] = 242;
// bram[30932] = 248;
// bram[30933] = 252;
// bram[30934] = 253;
// bram[30935] = 253;
// bram[30936] = 249;
// bram[30937] = 244;
// bram[30938] = 236;
// bram[30939] = 226;
// bram[30940] = 214;
// bram[30941] = 201;
// bram[30942] = 186;
// bram[30943] = 170;
// bram[30944] = 153;
// bram[30945] = 136;
// bram[30946] = 119;
// bram[30947] = 102;
// bram[30948] = 85;
// bram[30949] = 69;
// bram[30950] = 54;
// bram[30951] = 40;
// bram[30952] = 28;
// bram[30953] = 18;
// bram[30954] = 10;
// bram[30955] = 4;
// bram[30956] = 1;
// bram[30957] = 0;
// bram[30958] = 1;
// bram[30959] = 4;
// bram[30960] = 10;
// bram[30961] = 18;
// bram[30962] = 28;
// bram[30963] = 40;
// bram[30964] = 53;
// bram[30965] = 68;
// bram[30966] = 84;
// bram[30967] = 101;
// bram[30968] = 118;
// bram[30969] = 136;
// bram[30970] = 153;
// bram[30971] = 169;
// bram[30972] = 185;
// bram[30973] = 200;
// bram[30974] = 214;
// bram[30975] = 225;
// bram[30976] = 235;
// bram[30977] = 243;
// bram[30978] = 249;
// bram[30979] = 252;
// bram[30980] = 253;
// bram[30981] = 252;
// bram[30982] = 248;
// bram[30983] = 243;
// bram[30984] = 234;
// bram[30985] = 224;
// bram[30986] = 212;
// bram[30987] = 199;
// bram[30988] = 184;
// bram[30989] = 168;
// bram[30990] = 151;
// bram[30991] = 134;
// bram[30992] = 116;
// bram[30993] = 99;
// bram[30994] = 82;
// bram[30995] = 66;
// bram[30996] = 52;
// bram[30997] = 38;
// bram[30998] = 27;
// bram[30999] = 17;
// bram[31000] = 9;
// bram[31001] = 4;
// bram[31002] = 0;
// bram[31003] = 0;
// bram[31004] = 1;
// bram[31005] = 5;
// bram[31006] = 11;
// bram[31007] = 19;
// bram[31008] = 30;
// bram[31009] = 42;
// bram[31010] = 56;
// bram[31011] = 71;
// bram[31012] = 87;
// bram[31013] = 104;
// bram[31014] = 121;
// bram[31015] = 138;
// bram[31016] = 155;
// bram[31017] = 172;
// bram[31018] = 188;
// bram[31019] = 202;
// bram[31020] = 216;
// bram[31021] = 227;
// bram[31022] = 237;
// bram[31023] = 244;
// bram[31024] = 250;
// bram[31025] = 253;
// bram[31026] = 253;
// bram[31027] = 252;
// bram[31028] = 248;
// bram[31029] = 241;
// bram[31030] = 233;
// bram[31031] = 222;
// bram[31032] = 210;
// bram[31033] = 196;
// bram[31034] = 181;
// bram[31035] = 165;
// bram[31036] = 148;
// bram[31037] = 131;
// bram[31038] = 113;
// bram[31039] = 96;
// bram[31040] = 80;
// bram[31041] = 64;
// bram[31042] = 50;
// bram[31043] = 36;
// bram[31044] = 25;
// bram[31045] = 16;
// bram[31046] = 8;
// bram[31047] = 3;
// bram[31048] = 0;
// bram[31049] = 0;
// bram[31050] = 1;
// bram[31051] = 6;
// bram[31052] = 12;
// bram[31053] = 21;
// bram[31054] = 31;
// bram[31055] = 44;
// bram[31056] = 58;
// bram[31057] = 73;
// bram[31058] = 89;
// bram[31059] = 106;
// bram[31060] = 124;
// bram[31061] = 141;
// bram[31062] = 158;
// bram[31063] = 175;
// bram[31064] = 190;
// bram[31065] = 205;
// bram[31066] = 217;
// bram[31067] = 229;
// bram[31068] = 238;
// bram[31069] = 245;
// bram[31070] = 250;
// bram[31071] = 253;
// bram[31072] = 253;
// bram[31073] = 251;
// bram[31074] = 247;
// bram[31075] = 240;
// bram[31076] = 231;
// bram[31077] = 221;
// bram[31078] = 208;
// bram[31079] = 194;
// bram[31080] = 179;
// bram[31081] = 162;
// bram[31082] = 145;
// bram[31083] = 128;
// bram[31084] = 111;
// bram[31085] = 94;
// bram[31086] = 77;
// bram[31087] = 62;
// bram[31088] = 47;
// bram[31089] = 35;
// bram[31090] = 23;
// bram[31091] = 14;
// bram[31092] = 7;
// bram[31093] = 2;
// bram[31094] = 0;
// bram[31095] = 0;
// bram[31096] = 2;
// bram[31097] = 7;
// bram[31098] = 13;
// bram[31099] = 22;
// bram[31100] = 33;
// bram[31101] = 46;
// bram[31102] = 60;
// bram[31103] = 75;
// bram[31104] = 92;
// bram[31105] = 109;
// bram[31106] = 126;
// bram[31107] = 144;
// bram[31108] = 161;
// bram[31109] = 177;
// bram[31110] = 192;
// bram[31111] = 207;
// bram[31112] = 219;
// bram[31113] = 230;
// bram[31114] = 239;
// bram[31115] = 246;
// bram[31116] = 251;
// bram[31117] = 253;
// bram[31118] = 253;
// bram[31119] = 251;
// bram[31120] = 246;
// bram[31121] = 239;
// bram[31122] = 230;
// bram[31123] = 219;
// bram[31124] = 206;
// bram[31125] = 192;
// bram[31126] = 176;
// bram[31127] = 160;
// bram[31128] = 143;
// bram[31129] = 125;
// bram[31130] = 108;
// bram[31131] = 91;
// bram[31132] = 75;
// bram[31133] = 59;
// bram[31134] = 45;
// bram[31135] = 33;
// bram[31136] = 22;
// bram[31137] = 13;
// bram[31138] = 6;
// bram[31139] = 2;
// bram[31140] = 0;
// bram[31141] = 0;
// bram[31142] = 3;
// bram[31143] = 7;
// bram[31144] = 15;
// bram[31145] = 24;
// bram[31146] = 35;
// bram[31147] = 48;
// bram[31148] = 62;
// bram[31149] = 78;
// bram[31150] = 94;
// bram[31151] = 112;
// bram[31152] = 129;
// bram[31153] = 146;
// bram[31154] = 163;
// bram[31155] = 179;
// bram[31156] = 195;
// bram[31157] = 209;
// bram[31158] = 221;
// bram[31159] = 232;
// bram[31160] = 241;
// bram[31161] = 247;
// bram[31162] = 251;
// bram[31163] = 253;
// bram[31164] = 253;
// bram[31165] = 250;
// bram[31166] = 245;
// bram[31167] = 238;
// bram[31168] = 228;
// bram[31169] = 217;
// bram[31170] = 204;
// bram[31171] = 189;
// bram[31172] = 174;
// bram[31173] = 157;
// bram[31174] = 140;
// bram[31175] = 123;
// bram[31176] = 105;
// bram[31177] = 89;
// bram[31178] = 72;
// bram[31179] = 57;
// bram[31180] = 43;
// bram[31181] = 31;
// bram[31182] = 20;
// bram[31183] = 12;
// bram[31184] = 5;
// bram[31185] = 1;
// bram[31186] = 0;
// bram[31187] = 0;
// bram[31188] = 3;
// bram[31189] = 8;
// bram[31190] = 16;
// bram[31191] = 26;
// bram[31192] = 37;
// bram[31193] = 50;
// bram[31194] = 65;
// bram[31195] = 80;
// bram[31196] = 97;
// bram[31197] = 114;
// bram[31198] = 132;
// bram[31199] = 149;
// bram[31200] = 166;
// bram[31201] = 182;
// bram[31202] = 197;
// bram[31203] = 211;
// bram[31204] = 223;
// bram[31205] = 233;
// bram[31206] = 242;
// bram[31207] = 248;
// bram[31208] = 252;
// bram[31209] = 253;
// bram[31210] = 253;
// bram[31211] = 250;
// bram[31212] = 244;
// bram[31213] = 236;
// bram[31214] = 227;
// bram[31215] = 215;
// bram[31216] = 202;
// bram[31217] = 187;
// bram[31218] = 171;
// bram[31219] = 155;
// bram[31220] = 137;
// bram[31221] = 120;
// bram[31222] = 103;
// bram[31223] = 86;
// bram[31224] = 70;
// bram[31225] = 55;
// bram[31226] = 41;
// bram[31227] = 29;
// bram[31228] = 19;
// bram[31229] = 11;
// bram[31230] = 5;
// bram[31231] = 1;
// bram[31232] = 0;
// bram[31233] = 0;
// bram[31234] = 4;
// bram[31235] = 9;
// bram[31236] = 17;
// bram[31237] = 27;
// bram[31238] = 39;
// bram[31239] = 52;
// bram[31240] = 67;
// bram[31241] = 83;
// bram[31242] = 100;
// bram[31243] = 117;
// bram[31244] = 134;
// bram[31245] = 152;
// bram[31246] = 168;
// bram[31247] = 184;
// bram[31248] = 199;
// bram[31249] = 213;
// bram[31250] = 225;
// bram[31251] = 235;
// bram[31252] = 243;
// bram[31253] = 249;
// bram[31254] = 252;
// bram[31255] = 253;
// bram[31256] = 252;
// bram[31257] = 249;
// bram[31258] = 243;
// bram[31259] = 235;
// bram[31260] = 225;
// bram[31261] = 213;
// bram[31262] = 200;
// bram[31263] = 185;
// bram[31264] = 169;
// bram[31265] = 152;
// bram[31266] = 135;
// bram[31267] = 117;
// bram[31268] = 100;
// bram[31269] = 83;
// bram[31270] = 68;
// bram[31271] = 53;
// bram[31272] = 39;
// bram[31273] = 27;
// bram[31274] = 18;
// bram[31275] = 10;
// bram[31276] = 4;
// bram[31277] = 1;
// bram[31278] = 0;
// bram[31279] = 1;
// bram[31280] = 5;
// bram[31281] = 11;
// bram[31282] = 19;
// bram[31283] = 29;
// bram[31284] = 41;
// bram[31285] = 54;
// bram[31286] = 69;
// bram[31287] = 86;
// bram[31288] = 102;
// bram[31289] = 120;
// bram[31290] = 137;
// bram[31291] = 154;
// bram[31292] = 171;
// bram[31293] = 187;
// bram[31294] = 201;
// bram[31295] = 215;
// bram[31296] = 226;
// bram[31297] = 236;
// bram[31298] = 244;
// bram[31299] = 249;
// bram[31300] = 253;
// bram[31301] = 253;
// bram[31302] = 252;
// bram[31303] = 248;
// bram[31304] = 242;
// bram[31305] = 234;
// bram[31306] = 223;
// bram[31307] = 211;
// bram[31308] = 197;
// bram[31309] = 182;
// bram[31310] = 166;
// bram[31311] = 149;
// bram[31312] = 132;
// bram[31313] = 115;
// bram[31314] = 98;
// bram[31315] = 81;
// bram[31316] = 65;
// bram[31317] = 51;
// bram[31318] = 37;
// bram[31319] = 26;
// bram[31320] = 16;
// bram[31321] = 9;
// bram[31322] = 3;
// bram[31323] = 0;
// bram[31324] = 0;
// bram[31325] = 1;
// bram[31326] = 5;
// bram[31327] = 12;
// bram[31328] = 20;
// bram[31329] = 31;
// bram[31330] = 43;
// bram[31331] = 57;
// bram[31332] = 72;
// bram[31333] = 88;
// bram[31334] = 105;
// bram[31335] = 122;
// bram[31336] = 140;
// bram[31337] = 157;
// bram[31338] = 173;
// bram[31339] = 189;
// bram[31340] = 204;
// bram[31341] = 217;
// bram[31342] = 228;
// bram[31343] = 237;
// bram[31344] = 245;
// bram[31345] = 250;
// bram[31346] = 253;
// bram[31347] = 253;
// bram[31348] = 252;
// bram[31349] = 247;
// bram[31350] = 241;
// bram[31351] = 232;
// bram[31352] = 221;
// bram[31353] = 209;
// bram[31354] = 195;
// bram[31355] = 180;
// bram[31356] = 164;
// bram[31357] = 147;
// bram[31358] = 129;
// bram[31359] = 112;
// bram[31360] = 95;
// bram[31361] = 78;
// bram[31362] = 63;
// bram[31363] = 48;
// bram[31364] = 35;
// bram[31365] = 24;
// bram[31366] = 15;
// bram[31367] = 8;
// bram[31368] = 3;
// bram[31369] = 0;
// bram[31370] = 0;
// bram[31371] = 2;
// bram[31372] = 6;
// bram[31373] = 13;
// bram[31374] = 22;
// bram[31375] = 32;
// bram[31376] = 45;
// bram[31377] = 59;
// bram[31378] = 74;
// bram[31379] = 91;
// bram[31380] = 108;
// bram[31381] = 125;
// bram[31382] = 142;
// bram[31383] = 159;
// bram[31384] = 176;
// bram[31385] = 191;
// bram[31386] = 206;
// bram[31387] = 218;
// bram[31388] = 230;
// bram[31389] = 239;
// bram[31390] = 246;
// bram[31391] = 251;
// bram[31392] = 253;
// bram[31393] = 253;
// bram[31394] = 251;
// bram[31395] = 246;
// bram[31396] = 240;
// bram[31397] = 231;
// bram[31398] = 220;
// bram[31399] = 207;
// bram[31400] = 193;
// bram[31401] = 177;
// bram[31402] = 161;
// bram[31403] = 144;
// bram[31404] = 127;
// bram[31405] = 109;
// bram[31406] = 92;
// bram[31407] = 76;
// bram[31408] = 60;
// bram[31409] = 46;
// bram[31410] = 34;
// bram[31411] = 23;
// bram[31412] = 14;
// bram[31413] = 7;
// bram[31414] = 2;
// bram[31415] = 0;
// bram[31416] = 0;
// bram[31417] = 2;
// bram[31418] = 7;
// bram[31419] = 14;
// bram[31420] = 23;
// bram[31421] = 34;
// bram[31422] = 47;
// bram[31423] = 61;
// bram[31424] = 77;
// bram[31425] = 93;
// bram[31426] = 110;
// bram[31427] = 128;
// bram[31428] = 145;
// bram[31429] = 162;
// bram[31430] = 178;
// bram[31431] = 194;
// bram[31432] = 208;
// bram[31433] = 220;
// bram[31434] = 231;
// bram[31435] = 240;
// bram[31436] = 247;
// bram[31437] = 251;
// bram[31438] = 253;
// bram[31439] = 253;
// bram[31440] = 250;
// bram[31441] = 245;
// bram[31442] = 238;
// bram[31443] = 229;
// bram[31444] = 218;
// bram[31445] = 205;
// bram[31446] = 191;
// bram[31447] = 175;
// bram[31448] = 158;
// bram[31449] = 141;
// bram[31450] = 124;
// bram[31451] = 107;
// bram[31452] = 90;
// bram[31453] = 73;
// bram[31454] = 58;
// bram[31455] = 44;
// bram[31456] = 32;
// bram[31457] = 21;
// bram[31458] = 12;
// bram[31459] = 6;
// bram[31460] = 2;
// bram[31461] = 0;
// bram[31462] = 0;
// bram[31463] = 3;
// bram[31464] = 8;
// bram[31465] = 15;
// bram[31466] = 25;
// bram[31467] = 36;
// bram[31468] = 49;
// bram[31469] = 64;
// bram[31470] = 79;
// bram[31471] = 96;
// bram[31472] = 113;
// bram[31473] = 130;
// bram[31474] = 148;
// bram[31475] = 165;
// bram[31476] = 181;
// bram[31477] = 196;
// bram[31478] = 210;
// bram[31479] = 222;
// bram[31480] = 233;
// bram[31481] = 241;
// bram[31482] = 248;
// bram[31483] = 252;
// bram[31484] = 253;
// bram[31485] = 253;
// bram[31486] = 250;
// bram[31487] = 245;
// bram[31488] = 237;
// bram[31489] = 227;
// bram[31490] = 216;
// bram[31491] = 203;
// bram[31492] = 188;
// bram[31493] = 172;
// bram[31494] = 156;
// bram[31495] = 139;
// bram[31496] = 121;
// bram[31497] = 104;
// bram[31498] = 87;
// bram[31499] = 71;
// bram[31500] = 56;
// bram[31501] = 42;
// bram[31502] = 30;
// bram[31503] = 20;
// bram[31504] = 11;
// bram[31505] = 5;
// bram[31506] = 1;
// bram[31507] = 0;
// bram[31508] = 0;
// bram[31509] = 4;
// bram[31510] = 9;
// bram[31511] = 17;
// bram[31512] = 26;
// bram[31513] = 38;
// bram[31514] = 51;
// bram[31515] = 66;
// bram[31516] = 82;
// bram[31517] = 98;
// bram[31518] = 116;
// bram[31519] = 133;
// bram[31520] = 150;
// bram[31521] = 167;
// bram[31522] = 183;
// bram[31523] = 198;
// bram[31524] = 212;
// bram[31525] = 224;
// bram[31526] = 234;
// bram[31527] = 242;
// bram[31528] = 248;
// bram[31529] = 252;
// bram[31530] = 253;
// bram[31531] = 253;
// bram[31532] = 249;
// bram[31533] = 244;
// bram[31534] = 236;
// bram[31535] = 226;
// bram[31536] = 214;
// bram[31537] = 201;
// bram[31538] = 186;
// bram[31539] = 170;
// bram[31540] = 153;
// bram[31541] = 136;
// bram[31542] = 119;
// bram[31543] = 101;
// bram[31544] = 85;
// bram[31545] = 69;
// bram[31546] = 54;
// bram[31547] = 40;
// bram[31548] = 28;
// bram[31549] = 18;
// bram[31550] = 10;
// bram[31551] = 4;
// bram[31552] = 1;
// bram[31553] = 0;
// bram[31554] = 1;
// bram[31555] = 4;
// bram[31556] = 10;
// bram[31557] = 18;
// bram[31558] = 28;
// bram[31559] = 40;
// bram[31560] = 53;
// bram[31561] = 68;
// bram[31562] = 84;
// bram[31563] = 101;
// bram[31564] = 118;
// bram[31565] = 136;
// bram[31566] = 153;
// bram[31567] = 170;
// bram[31568] = 186;
// bram[31569] = 200;
// bram[31570] = 214;
// bram[31571] = 226;
// bram[31572] = 236;
// bram[31573] = 243;
// bram[31574] = 249;
// bram[31575] = 252;
// bram[31576] = 253;
// bram[31577] = 252;
// bram[31578] = 248;
// bram[31579] = 242;
// bram[31580] = 234;
// bram[31581] = 224;
// bram[31582] = 212;
// bram[31583] = 198;
// bram[31584] = 183;
// bram[31585] = 167;
// bram[31586] = 151;
// bram[31587] = 133;
// bram[31588] = 116;
// bram[31589] = 99;
// bram[31590] = 82;
// bram[31591] = 66;
// bram[31592] = 52;
// bram[31593] = 38;
// bram[31594] = 27;
// bram[31595] = 17;
// bram[31596] = 9;
// bram[31597] = 4;
// bram[31598] = 0;
// bram[31599] = 0;
// bram[31600] = 1;
// bram[31601] = 5;
// bram[31602] = 11;
// bram[31603] = 19;
// bram[31604] = 30;
// bram[31605] = 42;
// bram[31606] = 56;
// bram[31607] = 71;
// bram[31608] = 87;
// bram[31609] = 104;
// bram[31610] = 121;
// bram[31611] = 138;
// bram[31612] = 156;
// bram[31613] = 172;
// bram[31614] = 188;
// bram[31615] = 203;
// bram[31616] = 216;
// bram[31617] = 227;
// bram[31618] = 237;
// bram[31619] = 244;
// bram[31620] = 250;
// bram[31621] = 253;
// bram[31622] = 253;
// bram[31623] = 252;
// bram[31624] = 248;
// bram[31625] = 241;
// bram[31626] = 233;
// bram[31627] = 222;
// bram[31628] = 210;
// bram[31629] = 196;
// bram[31630] = 181;
// bram[31631] = 165;
// bram[31632] = 148;
// bram[31633] = 131;
// bram[31634] = 113;
// bram[31635] = 96;
// bram[31636] = 80;
// bram[31637] = 64;
// bram[31638] = 49;
// bram[31639] = 36;
// bram[31640] = 25;
// bram[31641] = 15;
// bram[31642] = 8;
// bram[31643] = 3;
// bram[31644] = 0;
// bram[31645] = 0;
// bram[31646] = 2;
// bram[31647] = 6;
// bram[31648] = 12;
// bram[31649] = 21;
// bram[31650] = 32;
// bram[31651] = 44;
// bram[31652] = 58;
// bram[31653] = 73;
// bram[31654] = 89;
// bram[31655] = 106;
// bram[31656] = 124;
// bram[31657] = 141;
// bram[31658] = 158;
// bram[31659] = 175;
// bram[31660] = 190;
// bram[31661] = 205;
// bram[31662] = 218;
// bram[31663] = 229;
// bram[31664] = 238;
// bram[31665] = 245;
// bram[31666] = 250;
// bram[31667] = 253;
// bram[31668] = 253;
// bram[31669] = 251;
// bram[31670] = 247;
// bram[31671] = 240;
// bram[31672] = 231;
// bram[31673] = 221;
// bram[31674] = 208;
// bram[31675] = 194;
// bram[31676] = 179;
// bram[31677] = 162;
// bram[31678] = 145;
// bram[31679] = 128;
// bram[31680] = 111;
// bram[31681] = 94;
// bram[31682] = 77;
// bram[31683] = 62;
// bram[31684] = 47;
// bram[31685] = 34;
// bram[31686] = 23;
// bram[31687] = 14;
// bram[31688] = 7;
// bram[31689] = 2;
// bram[31690] = 0;
// bram[31691] = 0;
// bram[31692] = 2;
// bram[31693] = 7;
// bram[31694] = 13;
// bram[31695] = 22;
// bram[31696] = 33;
// bram[31697] = 46;
// bram[31698] = 60;
// bram[31699] = 76;
// bram[31700] = 92;
// bram[31701] = 109;
// bram[31702] = 126;
// bram[31703] = 144;
// bram[31704] = 161;
// bram[31705] = 177;
// bram[31706] = 193;
// bram[31707] = 207;
// bram[31708] = 219;
// bram[31709] = 230;
// bram[31710] = 239;
// bram[31711] = 246;
// bram[31712] = 251;
// bram[31713] = 253;
// bram[31714] = 253;
// bram[31715] = 251;
// bram[31716] = 246;
// bram[31717] = 239;
// bram[31718] = 230;
// bram[31719] = 219;
// bram[31720] = 206;
// bram[31721] = 192;
// bram[31722] = 176;
// bram[31723] = 160;
// bram[31724] = 143;
// bram[31725] = 125;
// bram[31726] = 108;
// bram[31727] = 91;
// bram[31728] = 75;
// bram[31729] = 59;
// bram[31730] = 45;
// bram[31731] = 33;
// bram[31732] = 22;
// bram[31733] = 13;
// bram[31734] = 6;
// bram[31735] = 2;
// bram[31736] = 0;
// bram[31737] = 0;
// bram[31738] = 3;
// bram[31739] = 8;
// bram[31740] = 15;
// bram[31741] = 24;
// bram[31742] = 35;
// bram[31743] = 48;
// bram[31744] = 63;
// bram[31745] = 78;
// bram[31746] = 95;
// bram[31747] = 112;
// bram[31748] = 129;
// bram[31749] = 146;
// bram[31750] = 163;
// bram[31751] = 180;
// bram[31752] = 195;
// bram[31753] = 209;
// bram[31754] = 221;
// bram[31755] = 232;
// bram[31756] = 241;
// bram[31757] = 247;
// bram[31758] = 251;
// bram[31759] = 253;
// bram[31760] = 253;
// bram[31761] = 250;
// bram[31762] = 245;
// bram[31763] = 238;
// bram[31764] = 228;
// bram[31765] = 217;
// bram[31766] = 204;
// bram[31767] = 189;
// bram[31768] = 174;
// bram[31769] = 157;
// bram[31770] = 140;
// bram[31771] = 123;
// bram[31772] = 105;
// bram[31773] = 88;
// bram[31774] = 72;
// bram[31775] = 57;
// bram[31776] = 43;
// bram[31777] = 31;
// bram[31778] = 20;
// bram[31779] = 12;
// bram[31780] = 5;
// bram[31781] = 1;
// bram[31782] = 0;
// bram[31783] = 0;
// bram[31784] = 3;
// bram[31785] = 9;
// bram[31786] = 16;
// bram[31787] = 26;
// bram[31788] = 37;
// bram[31789] = 50;
// bram[31790] = 65;
// bram[31791] = 81;
// bram[31792] = 97;
// bram[31793] = 114;
// bram[31794] = 132;
// bram[31795] = 149;
// bram[31796] = 166;
// bram[31797] = 182;
// bram[31798] = 197;
// bram[31799] = 211;
// bram[31800] = 223;
// bram[31801] = 233;
// bram[31802] = 242;
// bram[31803] = 248;
// bram[31804] = 252;
// bram[31805] = 253;
// bram[31806] = 253;
// bram[31807] = 249;
// bram[31808] = 244;
// bram[31809] = 236;
// bram[31810] = 227;
// bram[31811] = 215;
// bram[31812] = 202;
// bram[31813] = 187;
// bram[31814] = 171;
// bram[31815] = 154;
// bram[31816] = 137;
// bram[31817] = 120;
// bram[31818] = 103;
// bram[31819] = 86;
// bram[31820] = 70;
// bram[31821] = 55;
// bram[31822] = 41;
// bram[31823] = 29;
// bram[31824] = 19;
// bram[31825] = 11;
// bram[31826] = 5;
// bram[31827] = 1;
// bram[31828] = 0;
// bram[31829] = 1;
// bram[31830] = 4;
// bram[31831] = 10;
// bram[31832] = 17;
// bram[31833] = 27;
// bram[31834] = 39;
// bram[31835] = 52;
// bram[31836] = 67;
// bram[31837] = 83;
// bram[31838] = 100;
// bram[31839] = 117;
// bram[31840] = 134;
// bram[31841] = 152;
// bram[31842] = 168;
// bram[31843] = 184;
// bram[31844] = 199;
// bram[31845] = 213;
// bram[31846] = 225;
// bram[31847] = 235;
// bram[31848] = 243;
// bram[31849] = 249;
// bram[31850] = 252;
// bram[31851] = 253;
// bram[31852] = 252;
// bram[31853] = 249;
// bram[31854] = 243;
// bram[31855] = 235;
// bram[31856] = 225;
// bram[31857] = 213;
// bram[31858] = 199;
// bram[31859] = 185;
// bram[31860] = 169;
// bram[31861] = 152;
// bram[31862] = 135;
// bram[31863] = 117;
// bram[31864] = 100;
// bram[31865] = 83;
// bram[31866] = 67;
// bram[31867] = 53;
// bram[31868] = 39;
// bram[31869] = 27;
// bram[31870] = 17;
// bram[31871] = 10;
// bram[31872] = 4;
// bram[31873] = 1;
// bram[31874] = 0;
// bram[31875] = 1;
// bram[31876] = 5;
// bram[31877] = 11;
// bram[31878] = 19;
// bram[31879] = 29;
// bram[31880] = 41;
// bram[31881] = 55;
// bram[31882] = 70;
// bram[31883] = 86;
// bram[31884] = 103;
// bram[31885] = 120;
// bram[31886] = 137;
// bram[31887] = 154;
// bram[31888] = 171;
// bram[31889] = 187;
// bram[31890] = 202;
// bram[31891] = 215;
// bram[31892] = 226;
// bram[31893] = 236;
// bram[31894] = 244;
// bram[31895] = 249;
// bram[31896] = 253;
// bram[31897] = 253;
// bram[31898] = 252;
// bram[31899] = 248;
// bram[31900] = 242;
// bram[31901] = 233;
// bram[31902] = 223;
// bram[31903] = 211;
// bram[31904] = 197;
// bram[31905] = 182;
// bram[31906] = 166;
// bram[31907] = 149;
// bram[31908] = 132;
// bram[31909] = 114;
// bram[31910] = 97;
// bram[31911] = 81;
// bram[31912] = 65;
// bram[31913] = 50;
// bram[31914] = 37;
// bram[31915] = 26;
// bram[31916] = 16;
// bram[31917] = 9;
// bram[31918] = 3;
// bram[31919] = 0;
// bram[31920] = 0;
// bram[31921] = 1;
// bram[31922] = 5;
// bram[31923] = 12;
// bram[31924] = 20;
// bram[31925] = 31;
// bram[31926] = 43;
// bram[31927] = 57;
// bram[31928] = 72;
// bram[31929] = 88;
// bram[31930] = 105;
// bram[31931] = 122;
// bram[31932] = 140;
// bram[31933] = 157;
// bram[31934] = 174;
// bram[31935] = 189;
// bram[31936] = 204;
// bram[31937] = 217;
// bram[31938] = 228;
// bram[31939] = 238;
// bram[31940] = 245;
// bram[31941] = 250;
// bram[31942] = 253;
// bram[31943] = 253;
// bram[31944] = 251;
// bram[31945] = 247;
// bram[31946] = 241;
// bram[31947] = 232;
// bram[31948] = 221;
// bram[31949] = 209;
// bram[31950] = 195;
// bram[31951] = 180;
// bram[31952] = 163;
// bram[31953] = 147;
// bram[31954] = 129;
// bram[31955] = 112;
// bram[31956] = 95;
// bram[31957] = 78;
// bram[31958] = 63;
// bram[31959] = 48;
// bram[31960] = 35;
// bram[31961] = 24;
// bram[31962] = 15;
// bram[31963] = 8;
// bram[31964] = 3;
// bram[31965] = 0;
// bram[31966] = 0;
// bram[31967] = 2;
// bram[31968] = 6;
// bram[31969] = 13;
// bram[31970] = 22;
// bram[31971] = 33;
// bram[31972] = 45;
// bram[31973] = 59;
// bram[31974] = 75;
// bram[31975] = 91;
// bram[31976] = 108;
// bram[31977] = 125;
// bram[31978] = 143;
// bram[31979] = 160;
// bram[31980] = 176;
// bram[31981] = 192;
// bram[31982] = 206;
// bram[31983] = 219;
// bram[31984] = 230;
// bram[31985] = 239;
// bram[31986] = 246;
// bram[31987] = 251;
// bram[31988] = 253;
// bram[31989] = 253;
// bram[31990] = 251;
// bram[31991] = 246;
// bram[31992] = 239;
// bram[31993] = 230;
// bram[31994] = 220;
// bram[31995] = 207;
// bram[31996] = 193;
// bram[31997] = 177;
// bram[31998] = 161;
// bram[31999] = 144;
// bram[32000] = 127;
// bram[32001] = 146;
// bram[32002] = 165;
// bram[32003] = 183;
// bram[32004] = 200;
// bram[32005] = 215;
// bram[32006] = 228;
// bram[32007] = 238;
// bram[32008] = 246;
// bram[32009] = 251;
// bram[32010] = 253;
// bram[32011] = 253;
// bram[32012] = 249;
// bram[32013] = 242;
// bram[32014] = 232;
// bram[32015] = 220;
// bram[32016] = 206;
// bram[32017] = 190;
// bram[32018] = 173;
// bram[32019] = 154;
// bram[32020] = 134;
// bram[32021] = 115;
// bram[32022] = 96;
// bram[32023] = 77;
// bram[32024] = 60;
// bram[32025] = 44;
// bram[32026] = 30;
// bram[32027] = 19;
// bram[32028] = 10;
// bram[32029] = 3;
// bram[32030] = 0;
// bram[32031] = 0;
// bram[32032] = 2;
// bram[32033] = 8;
// bram[32034] = 16;
// bram[32035] = 27;
// bram[32036] = 41;
// bram[32037] = 56;
// bram[32038] = 73;
// bram[32039] = 91;
// bram[32040] = 111;
// bram[32041] = 130;
// bram[32042] = 150;
// bram[32043] = 168;
// bram[32044] = 186;
// bram[32045] = 203;
// bram[32046] = 217;
// bram[32047] = 230;
// bram[32048] = 240;
// bram[32049] = 247;
// bram[32050] = 252;
// bram[32051] = 253;
// bram[32052] = 252;
// bram[32053] = 248;
// bram[32054] = 240;
// bram[32055] = 230;
// bram[32056] = 218;
// bram[32057] = 203;
// bram[32058] = 187;
// bram[32059] = 169;
// bram[32060] = 150;
// bram[32061] = 131;
// bram[32062] = 111;
// bram[32063] = 92;
// bram[32064] = 74;
// bram[32065] = 57;
// bram[32066] = 41;
// bram[32067] = 28;
// bram[32068] = 17;
// bram[32069] = 8;
// bram[32070] = 3;
// bram[32071] = 0;
// bram[32072] = 0;
// bram[32073] = 3;
// bram[32074] = 9;
// bram[32075] = 18;
// bram[32076] = 30;
// bram[32077] = 43;
// bram[32078] = 59;
// bram[32079] = 76;
// bram[32080] = 95;
// bram[32081] = 114;
// bram[32082] = 134;
// bram[32083] = 153;
// bram[32084] = 172;
// bram[32085] = 189;
// bram[32086] = 206;
// bram[32087] = 220;
// bram[32088] = 232;
// bram[32089] = 242;
// bram[32090] = 248;
// bram[32091] = 252;
// bram[32092] = 253;
// bram[32093] = 251;
// bram[32094] = 247;
// bram[32095] = 239;
// bram[32096] = 228;
// bram[32097] = 215;
// bram[32098] = 201;
// bram[32099] = 184;
// bram[32100] = 166;
// bram[32101] = 147;
// bram[32102] = 127;
// bram[32103] = 108;
// bram[32104] = 89;
// bram[32105] = 71;
// bram[32106] = 54;
// bram[32107] = 39;
// bram[32108] = 26;
// bram[32109] = 15;
// bram[32110] = 7;
// bram[32111] = 2;
// bram[32112] = 0;
// bram[32113] = 0;
// bram[32114] = 4;
// bram[32115] = 11;
// bram[32116] = 20;
// bram[32117] = 32;
// bram[32118] = 46;
// bram[32119] = 62;
// bram[32120] = 80;
// bram[32121] = 98;
// bram[32122] = 118;
// bram[32123] = 137;
// bram[32124] = 157;
// bram[32125] = 175;
// bram[32126] = 193;
// bram[32127] = 208;
// bram[32128] = 222;
// bram[32129] = 234;
// bram[32130] = 243;
// bram[32131] = 249;
// bram[32132] = 253;
// bram[32133] = 253;
// bram[32134] = 251;
// bram[32135] = 245;
// bram[32136] = 237;
// bram[32137] = 226;
// bram[32138] = 213;
// bram[32139] = 198;
// bram[32140] = 181;
// bram[32141] = 162;
// bram[32142] = 143;
// bram[32143] = 124;
// bram[32144] = 104;
// bram[32145] = 85;
// bram[32146] = 67;
// bram[32147] = 51;
// bram[32148] = 36;
// bram[32149] = 24;
// bram[32150] = 13;
// bram[32151] = 6;
// bram[32152] = 1;
// bram[32153] = 0;
// bram[32154] = 1;
// bram[32155] = 5;
// bram[32156] = 12;
// bram[32157] = 22;
// bram[32158] = 34;
// bram[32159] = 49;
// bram[32160] = 65;
// bram[32161] = 83;
// bram[32162] = 102;
// bram[32163] = 121;
// bram[32164] = 141;
// bram[32165] = 160;
// bram[32166] = 178;
// bram[32167] = 196;
// bram[32168] = 211;
// bram[32169] = 225;
// bram[32170] = 236;
// bram[32171] = 244;
// bram[32172] = 250;
// bram[32173] = 253;
// bram[32174] = 253;
// bram[32175] = 250;
// bram[32176] = 244;
// bram[32177] = 235;
// bram[32178] = 224;
// bram[32179] = 210;
// bram[32180] = 195;
// bram[32181] = 177;
// bram[32182] = 159;
// bram[32183] = 140;
// bram[32184] = 120;
// bram[32185] = 101;
// bram[32186] = 82;
// bram[32187] = 64;
// bram[32188] = 48;
// bram[32189] = 34;
// bram[32190] = 21;
// bram[32191] = 12;
// bram[32192] = 5;
// bram[32193] = 1;
// bram[32194] = 0;
// bram[32195] = 1;
// bram[32196] = 6;
// bram[32197] = 14;
// bram[32198] = 24;
// bram[32199] = 37;
// bram[32200] = 52;
// bram[32201] = 68;
// bram[32202] = 86;
// bram[32203] = 105;
// bram[32204] = 125;
// bram[32205] = 144;
// bram[32206] = 163;
// bram[32207] = 182;
// bram[32208] = 199;
// bram[32209] = 214;
// bram[32210] = 227;
// bram[32211] = 238;
// bram[32212] = 246;
// bram[32213] = 251;
// bram[32214] = 253;
// bram[32215] = 253;
// bram[32216] = 249;
// bram[32217] = 243;
// bram[32218] = 233;
// bram[32219] = 221;
// bram[32220] = 207;
// bram[32221] = 191;
// bram[32222] = 174;
// bram[32223] = 155;
// bram[32224] = 136;
// bram[32225] = 117;
// bram[32226] = 97;
// bram[32227] = 79;
// bram[32228] = 61;
// bram[32229] = 45;
// bram[32230] = 31;
// bram[32231] = 19;
// bram[32232] = 10;
// bram[32233] = 4;
// bram[32234] = 0;
// bram[32235] = 0;
// bram[32236] = 2;
// bram[32237] = 7;
// bram[32238] = 16;
// bram[32239] = 26;
// bram[32240] = 40;
// bram[32241] = 55;
// bram[32242] = 72;
// bram[32243] = 90;
// bram[32244] = 109;
// bram[32245] = 128;
// bram[32246] = 148;
// bram[32247] = 167;
// bram[32248] = 185;
// bram[32249] = 201;
// bram[32250] = 216;
// bram[32251] = 229;
// bram[32252] = 239;
// bram[32253] = 247;
// bram[32254] = 252;
// bram[32255] = 253;
// bram[32256] = 252;
// bram[32257] = 248;
// bram[32258] = 241;
// bram[32259] = 231;
// bram[32260] = 219;
// bram[32261] = 205;
// bram[32262] = 188;
// bram[32263] = 171;
// bram[32264] = 152;
// bram[32265] = 132;
// bram[32266] = 113;
// bram[32267] = 94;
// bram[32268] = 75;
// bram[32269] = 58;
// bram[32270] = 43;
// bram[32271] = 29;
// bram[32272] = 18;
// bram[32273] = 9;
// bram[32274] = 3;
// bram[32275] = 0;
// bram[32276] = 0;
// bram[32277] = 3;
// bram[32278] = 9;
// bram[32279] = 17;
// bram[32280] = 29;
// bram[32281] = 42;
// bram[32282] = 58;
// bram[32283] = 75;
// bram[32284] = 93;
// bram[32285] = 113;
// bram[32286] = 132;
// bram[32287] = 151;
// bram[32288] = 170;
// bram[32289] = 188;
// bram[32290] = 204;
// bram[32291] = 219;
// bram[32292] = 231;
// bram[32293] = 241;
// bram[32294] = 248;
// bram[32295] = 252;
// bram[32296] = 253;
// bram[32297] = 252;
// bram[32298] = 247;
// bram[32299] = 239;
// bram[32300] = 229;
// bram[32301] = 217;
// bram[32302] = 202;
// bram[32303] = 185;
// bram[32304] = 167;
// bram[32305] = 148;
// bram[32306] = 129;
// bram[32307] = 109;
// bram[32308] = 90;
// bram[32309] = 72;
// bram[32310] = 55;
// bram[32311] = 40;
// bram[32312] = 27;
// bram[32313] = 16;
// bram[32314] = 8;
// bram[32315] = 2;
// bram[32316] = 0;
// bram[32317] = 0;
// bram[32318] = 4;
// bram[32319] = 10;
// bram[32320] = 19;
// bram[32321] = 31;
// bram[32322] = 45;
// bram[32323] = 61;
// bram[32324] = 78;
// bram[32325] = 97;
// bram[32326] = 116;
// bram[32327] = 136;
// bram[32328] = 155;
// bram[32329] = 174;
// bram[32330] = 191;
// bram[32331] = 207;
// bram[32332] = 221;
// bram[32333] = 233;
// bram[32334] = 242;
// bram[32335] = 249;
// bram[32336] = 253;
// bram[32337] = 253;
// bram[32338] = 251;
// bram[32339] = 246;
// bram[32340] = 238;
// bram[32341] = 227;
// bram[32342] = 214;
// bram[32343] = 199;
// bram[32344] = 182;
// bram[32345] = 164;
// bram[32346] = 145;
// bram[32347] = 125;
// bram[32348] = 106;
// bram[32349] = 87;
// bram[32350] = 69;
// bram[32351] = 52;
// bram[32352] = 37;
// bram[32353] = 24;
// bram[32354] = 14;
// bram[32355] = 6;
// bram[32356] = 1;
// bram[32357] = 0;
// bram[32358] = 1;
// bram[32359] = 5;
// bram[32360] = 12;
// bram[32361] = 21;
// bram[32362] = 33;
// bram[32363] = 48;
// bram[32364] = 64;
// bram[32365] = 82;
// bram[32366] = 100;
// bram[32367] = 120;
// bram[32368] = 139;
// bram[32369] = 158;
// bram[32370] = 177;
// bram[32371] = 194;
// bram[32372] = 210;
// bram[32373] = 224;
// bram[32374] = 235;
// bram[32375] = 244;
// bram[32376] = 250;
// bram[32377] = 253;
// bram[32378] = 253;
// bram[32379] = 250;
// bram[32380] = 245;
// bram[32381] = 236;
// bram[32382] = 225;
// bram[32383] = 211;
// bram[32384] = 196;
// bram[32385] = 179;
// bram[32386] = 160;
// bram[32387] = 141;
// bram[32388] = 122;
// bram[32389] = 102;
// bram[32390] = 83;
// bram[32391] = 66;
// bram[32392] = 49;
// bram[32393] = 35;
// bram[32394] = 22;
// bram[32395] = 12;
// bram[32396] = 5;
// bram[32397] = 1;
// bram[32398] = 0;
// bram[32399] = 1;
// bram[32400] = 6;
// bram[32401] = 13;
// bram[32402] = 23;
// bram[32403] = 36;
// bram[32404] = 51;
// bram[32405] = 67;
// bram[32406] = 85;
// bram[32407] = 104;
// bram[32408] = 123;
// bram[32409] = 143;
// bram[32410] = 162;
// bram[32411] = 180;
// bram[32412] = 197;
// bram[32413] = 213;
// bram[32414] = 226;
// bram[32415] = 237;
// bram[32416] = 245;
// bram[32417] = 251;
// bram[32418] = 253;
// bram[32419] = 253;
// bram[32420] = 250;
// bram[32421] = 243;
// bram[32422] = 234;
// bram[32423] = 223;
// bram[32424] = 209;
// bram[32425] = 193;
// bram[32426] = 175;
// bram[32427] = 157;
// bram[32428] = 138;
// bram[32429] = 118;
// bram[32430] = 99;
// bram[32431] = 80;
// bram[32432] = 63;
// bram[32433] = 46;
// bram[32434] = 32;
// bram[32435] = 20;
// bram[32436] = 11;
// bram[32437] = 4;
// bram[32438] = 0;
// bram[32439] = 0;
// bram[32440] = 2;
// bram[32441] = 7;
// bram[32442] = 15;
// bram[32443] = 25;
// bram[32444] = 38;
// bram[32445] = 53;
// bram[32446] = 70;
// bram[32447] = 88;
// bram[32448] = 107;
// bram[32449] = 127;
// bram[32450] = 146;
// bram[32451] = 165;
// bram[32452] = 183;
// bram[32453] = 200;
// bram[32454] = 215;
// bram[32455] = 228;
// bram[32456] = 239;
// bram[32457] = 246;
// bram[32458] = 251;
// bram[32459] = 253;
// bram[32460] = 252;
// bram[32461] = 249;
// bram[32462] = 242;
// bram[32463] = 232;
// bram[32464] = 220;
// bram[32465] = 206;
// bram[32466] = 190;
// bram[32467] = 172;
// bram[32468] = 153;
// bram[32469] = 134;
// bram[32470] = 115;
// bram[32471] = 95;
// bram[32472] = 77;
// bram[32473] = 59;
// bram[32474] = 44;
// bram[32475] = 30;
// bram[32476] = 18;
// bram[32477] = 9;
// bram[32478] = 3;
// bram[32479] = 0;
// bram[32480] = 0;
// bram[32481] = 2;
// bram[32482] = 8;
// bram[32483] = 17;
// bram[32484] = 28;
// bram[32485] = 41;
// bram[32486] = 56;
// bram[32487] = 74;
// bram[32488] = 92;
// bram[32489] = 111;
// bram[32490] = 130;
// bram[32491] = 150;
// bram[32492] = 169;
// bram[32493] = 187;
// bram[32494] = 203;
// bram[32495] = 218;
// bram[32496] = 230;
// bram[32497] = 240;
// bram[32498] = 248;
// bram[32499] = 252;
// bram[32500] = 254;
// bram[32501] = 252;
// bram[32502] = 248;
// bram[32503] = 240;
// bram[32504] = 230;
// bram[32505] = 218;
// bram[32506] = 203;
// bram[32507] = 187;
// bram[32508] = 169;
// bram[32509] = 150;
// bram[32510] = 130;
// bram[32511] = 111;
// bram[32512] = 92;
// bram[32513] = 74;
// bram[32514] = 56;
// bram[32515] = 41;
// bram[32516] = 28;
// bram[32517] = 17;
// bram[32518] = 8;
// bram[32519] = 2;
// bram[32520] = 0;
// bram[32521] = 0;
// bram[32522] = 3;
// bram[32523] = 9;
// bram[32524] = 18;
// bram[32525] = 30;
// bram[32526] = 44;
// bram[32527] = 59;
// bram[32528] = 77;
// bram[32529] = 95;
// bram[32530] = 115;
// bram[32531] = 134;
// bram[32532] = 153;
// bram[32533] = 172;
// bram[32534] = 190;
// bram[32535] = 206;
// bram[32536] = 220;
// bram[32537] = 232;
// bram[32538] = 242;
// bram[32539] = 249;
// bram[32540] = 252;
// bram[32541] = 253;
// bram[32542] = 251;
// bram[32543] = 246;
// bram[32544] = 239;
// bram[32545] = 228;
// bram[32546] = 215;
// bram[32547] = 200;
// bram[32548] = 183;
// bram[32549] = 165;
// bram[32550] = 146;
// bram[32551] = 127;
// bram[32552] = 107;
// bram[32553] = 88;
// bram[32554] = 70;
// bram[32555] = 53;
// bram[32556] = 38;
// bram[32557] = 25;
// bram[32558] = 15;
// bram[32559] = 7;
// bram[32560] = 2;
// bram[32561] = 0;
// bram[32562] = 0;
// bram[32563] = 4;
// bram[32564] = 11;
// bram[32565] = 20;
// bram[32566] = 32;
// bram[32567] = 46;
// bram[32568] = 63;
// bram[32569] = 80;
// bram[32570] = 99;
// bram[32571] = 118;
// bram[32572] = 138;
// bram[32573] = 157;
// bram[32574] = 175;
// bram[32575] = 193;
// bram[32576] = 209;
// bram[32577] = 223;
// bram[32578] = 234;
// bram[32579] = 243;
// bram[32580] = 250;
// bram[32581] = 253;
// bram[32582] = 253;
// bram[32583] = 251;
// bram[32584] = 245;
// bram[32585] = 237;
// bram[32586] = 226;
// bram[32587] = 213;
// bram[32588] = 197;
// bram[32589] = 180;
// bram[32590] = 162;
// bram[32591] = 143;
// bram[32592] = 123;
// bram[32593] = 104;
// bram[32594] = 85;
// bram[32595] = 67;
// bram[32596] = 51;
// bram[32597] = 36;
// bram[32598] = 23;
// bram[32599] = 13;
// bram[32600] = 6;
// bram[32601] = 1;
// bram[32602] = 0;
// bram[32603] = 1;
// bram[32604] = 5;
// bram[32605] = 12;
// bram[32606] = 22;
// bram[32607] = 35;
// bram[32608] = 49;
// bram[32609] = 66;
// bram[32610] = 83;
// bram[32611] = 102;
// bram[32612] = 122;
// bram[32613] = 141;
// bram[32614] = 160;
// bram[32615] = 179;
// bram[32616] = 196;
// bram[32617] = 211;
// bram[32618] = 225;
// bram[32619] = 236;
// bram[32620] = 245;
// bram[32621] = 250;
// bram[32622] = 253;
// bram[32623] = 253;
// bram[32624] = 250;
// bram[32625] = 244;
// bram[32626] = 235;
// bram[32627] = 224;
// bram[32628] = 210;
// bram[32629] = 194;
// bram[32630] = 177;
// bram[32631] = 158;
// bram[32632] = 139;
// bram[32633] = 120;
// bram[32634] = 100;
// bram[32635] = 82;
// bram[32636] = 64;
// bram[32637] = 48;
// bram[32638] = 33;
// bram[32639] = 21;
// bram[32640] = 12;
// bram[32641] = 5;
// bram[32642] = 1;
// bram[32643] = 0;
// bram[32644] = 1;
// bram[32645] = 6;
// bram[32646] = 14;
// bram[32647] = 24;
// bram[32648] = 37;
// bram[32649] = 52;
// bram[32650] = 69;
// bram[32651] = 87;
// bram[32652] = 106;
// bram[32653] = 125;
// bram[32654] = 145;
// bram[32655] = 164;
// bram[32656] = 182;
// bram[32657] = 199;
// bram[32658] = 214;
// bram[32659] = 227;
// bram[32660] = 238;
// bram[32661] = 246;
// bram[32662] = 251;
// bram[32663] = 253;
// bram[32664] = 253;
// bram[32665] = 249;
// bram[32666] = 242;
// bram[32667] = 233;
// bram[32668] = 221;
// bram[32669] = 207;
// bram[32670] = 191;
// bram[32671] = 174;
// bram[32672] = 155;
// bram[32673] = 136;
// bram[32674] = 116;
// bram[32675] = 97;
// bram[32676] = 78;
// bram[32677] = 61;
// bram[32678] = 45;
// bram[32679] = 31;
// bram[32680] = 19;
// bram[32681] = 10;
// bram[32682] = 4;
// bram[32683] = 0;
// bram[32684] = 0;
// bram[32685] = 2;
// bram[32686] = 8;
// bram[32687] = 16;
// bram[32688] = 27;
// bram[32689] = 40;
// bram[32690] = 55;
// bram[32691] = 72;
// bram[32692] = 90;
// bram[32693] = 109;
// bram[32694] = 129;
// bram[32695] = 148;
// bram[32696] = 167;
// bram[32697] = 185;
// bram[32698] = 202;
// bram[32699] = 217;
// bram[32700] = 229;
// bram[32701] = 239;
// bram[32702] = 247;
// bram[32703] = 252;
// bram[32704] = 253;
// bram[32705] = 252;
// bram[32706] = 248;
// bram[32707] = 241;
// bram[32708] = 231;
// bram[32709] = 219;
// bram[32710] = 204;
// bram[32711] = 188;
// bram[32712] = 170;
// bram[32713] = 151;
// bram[32714] = 132;
// bram[32715] = 113;
// bram[32716] = 93;
// bram[32717] = 75;
// bram[32718] = 58;
// bram[32719] = 42;
// bram[32720] = 29;
// bram[32721] = 17;
// bram[32722] = 9;
// bram[32723] = 3;
// bram[32724] = 0;
// bram[32725] = 0;
// bram[32726] = 3;
// bram[32727] = 9;
// bram[32728] = 18;
// bram[32729] = 29;
// bram[32730] = 43;
// bram[32731] = 58;
// bram[32732] = 75;
// bram[32733] = 94;
// bram[32734] = 113;
// bram[32735] = 132;
// bram[32736] = 152;
// bram[32737] = 171;
// bram[32738] = 188;
// bram[32739] = 205;
// bram[32740] = 219;
// bram[32741] = 231;
// bram[32742] = 241;
// bram[32743] = 248;
// bram[32744] = 252;
// bram[32745] = 253;
// bram[32746] = 252;
// bram[32747] = 247;
// bram[32748] = 239;
// bram[32749] = 229;
// bram[32750] = 216;
// bram[32751] = 201;
// bram[32752] = 185;
// bram[32753] = 167;
// bram[32754] = 148;
// bram[32755] = 128;
// bram[32756] = 109;
// bram[32757] = 90;
// bram[32758] = 72;
// bram[32759] = 55;
// bram[32760] = 40;
// bram[32761] = 26;
// bram[32762] = 16;
// bram[32763] = 7;
// bram[32764] = 2;
// bram[32765] = 0;
// bram[32766] = 0;
// bram[32767] = 4;
// bram[32768] = 10;
// bram[32769] = 19;
// bram[32770] = 31;
// bram[32771] = 45;
// bram[32772] = 61;
// bram[32773] = 79;
// bram[32774] = 97;
// bram[32775] = 117;
// bram[32776] = 136;
// bram[32777] = 155;
// bram[32778] = 174;
// bram[32779] = 191;
// bram[32780] = 207;
// bram[32781] = 221;
// bram[32782] = 233;
// bram[32783] = 243;
// bram[32784] = 249;
// bram[32785] = 253;
// bram[32786] = 253;
// bram[32787] = 251;
// bram[32788] = 246;
// bram[32789] = 238;
// bram[32790] = 227;
// bram[32791] = 214;
// bram[32792] = 199;
// bram[32793] = 182;
// bram[32794] = 163;
// bram[32795] = 144;
// bram[32796] = 125;
// bram[32797] = 105;
// bram[32798] = 86;
// bram[32799] = 68;
// bram[32800] = 52;
// bram[32801] = 37;
// bram[32802] = 24;
// bram[32803] = 14;
// bram[32804] = 6;
// bram[32805] = 1;
// bram[32806] = 0;
// bram[32807] = 1;
// bram[32808] = 5;
// bram[32809] = 12;
// bram[32810] = 21;
// bram[32811] = 34;
// bram[32812] = 48;
// bram[32813] = 64;
// bram[32814] = 82;
// bram[32815] = 101;
// bram[32816] = 120;
// bram[32817] = 140;
// bram[32818] = 159;
// bram[32819] = 177;
// bram[32820] = 195;
// bram[32821] = 210;
// bram[32822] = 224;
// bram[32823] = 235;
// bram[32824] = 244;
// bram[32825] = 250;
// bram[32826] = 253;
// bram[32827] = 253;
// bram[32828] = 250;
// bram[32829] = 244;
// bram[32830] = 236;
// bram[32831] = 225;
// bram[32832] = 211;
// bram[32833] = 196;
// bram[32834] = 178;
// bram[32835] = 160;
// bram[32836] = 141;
// bram[32837] = 121;
// bram[32838] = 102;
// bram[32839] = 83;
// bram[32840] = 65;
// bram[32841] = 49;
// bram[32842] = 34;
// bram[32843] = 22;
// bram[32844] = 12;
// bram[32845] = 5;
// bram[32846] = 1;
// bram[32847] = 0;
// bram[32848] = 1;
// bram[32849] = 6;
// bram[32850] = 13;
// bram[32851] = 24;
// bram[32852] = 36;
// bram[32853] = 51;
// bram[32854] = 67;
// bram[32855] = 85;
// bram[32856] = 104;
// bram[32857] = 124;
// bram[32858] = 143;
// bram[32859] = 162;
// bram[32860] = 181;
// bram[32861] = 198;
// bram[32862] = 213;
// bram[32863] = 226;
// bram[32864] = 237;
// bram[32865] = 245;
// bram[32866] = 251;
// bram[32867] = 253;
// bram[32868] = 253;
// bram[32869] = 249;
// bram[32870] = 243;
// bram[32871] = 234;
// bram[32872] = 222;
// bram[32873] = 208;
// bram[32874] = 193;
// bram[32875] = 175;
// bram[32876] = 157;
// bram[32877] = 137;
// bram[32878] = 118;
// bram[32879] = 98;
// bram[32880] = 80;
// bram[32881] = 62;
// bram[32882] = 46;
// bram[32883] = 32;
// bram[32884] = 20;
// bram[32885] = 11;
// bram[32886] = 4;
// bram[32887] = 0;
// bram[32888] = 0;
// bram[32889] = 2;
// bram[32890] = 7;
// bram[32891] = 15;
// bram[32892] = 26;
// bram[32893] = 39;
// bram[32894] = 54;
// bram[32895] = 71;
// bram[32896] = 89;
// bram[32897] = 108;
// bram[32898] = 127;
// bram[32899] = 147;
// bram[32900] = 166;
// bram[32901] = 184;
// bram[32902] = 201;
// bram[32903] = 215;
// bram[32904] = 228;
// bram[32905] = 239;
// bram[32906] = 247;
// bram[32907] = 251;
// bram[32908] = 253;
// bram[32909] = 252;
// bram[32910] = 248;
// bram[32911] = 242;
// bram[32912] = 232;
// bram[32913] = 220;
// bram[32914] = 206;
// bram[32915] = 189;
// bram[32916] = 172;
// bram[32917] = 153;
// bram[32918] = 134;
// bram[32919] = 114;
// bram[32920] = 95;
// bram[32921] = 76;
// bram[32922] = 59;
// bram[32923] = 43;
// bram[32924] = 30;
// bram[32925] = 18;
// bram[32926] = 9;
// bram[32927] = 3;
// bram[32928] = 0;
// bram[32929] = 0;
// bram[32930] = 3;
// bram[32931] = 8;
// bram[32932] = 17;
// bram[32933] = 28;
// bram[32934] = 41;
// bram[32935] = 57;
// bram[32936] = 74;
// bram[32937] = 92;
// bram[32938] = 111;
// bram[32939] = 131;
// bram[32940] = 150;
// bram[32941] = 169;
// bram[32942] = 187;
// bram[32943] = 203;
// bram[32944] = 218;
// bram[32945] = 230;
// bram[32946] = 240;
// bram[32947] = 248;
// bram[32948] = 252;
// bram[32949] = 253;
// bram[32950] = 252;
// bram[32951] = 247;
// bram[32952] = 240;
// bram[32953] = 230;
// bram[32954] = 217;
// bram[32955] = 203;
// bram[32956] = 186;
// bram[32957] = 168;
// bram[32958] = 150;
// bram[32959] = 130;
// bram[32960] = 111;
// bram[32961] = 91;
// bram[32962] = 73;
// bram[32963] = 56;
// bram[32964] = 41;
// bram[32965] = 27;
// bram[32966] = 16;
// bram[32967] = 8;
// bram[32968] = 2;
// bram[32969] = 0;
// bram[32970] = 0;
// bram[32971] = 3;
// bram[32972] = 10;
// bram[32973] = 19;
// bram[32974] = 30;
// bram[32975] = 44;
// bram[32976] = 60;
// bram[32977] = 77;
// bram[32978] = 96;
// bram[32979] = 115;
// bram[32980] = 134;
// bram[32981] = 154;
// bram[32982] = 173;
// bram[32983] = 190;
// bram[32984] = 206;
// bram[32985] = 220;
// bram[32986] = 232;
// bram[32987] = 242;
// bram[32988] = 249;
// bram[32989] = 253;
// bram[32990] = 253;
// bram[32991] = 251;
// bram[32992] = 246;
// bram[32993] = 238;
// bram[32994] = 228;
// bram[32995] = 215;
// bram[32996] = 200;
// bram[32997] = 183;
// bram[32998] = 165;
// bram[32999] = 146;
// bram[33000] = 127;
// bram[33001] = 107;
// bram[33002] = 88;
// bram[33003] = 70;
// bram[33004] = 53;
// bram[33005] = 38;
// bram[33006] = 25;
// bram[33007] = 15;
// bram[33008] = 7;
// bram[33009] = 2;
// bram[33010] = 0;
// bram[33011] = 0;
// bram[33012] = 4;
// bram[33013] = 11;
// bram[33014] = 21;
// bram[33015] = 33;
// bram[33016] = 47;
// bram[33017] = 63;
// bram[33018] = 80;
// bram[33019] = 99;
// bram[33020] = 119;
// bram[33021] = 138;
// bram[33022] = 157;
// bram[33023] = 176;
// bram[33024] = 193;
// bram[33025] = 209;
// bram[33026] = 223;
// bram[33027] = 234;
// bram[33028] = 243;
// bram[33029] = 250;
// bram[33030] = 253;
// bram[33031] = 253;
// bram[33032] = 251;
// bram[33033] = 245;
// bram[33034] = 237;
// bram[33035] = 226;
// bram[33036] = 212;
// bram[33037] = 197;
// bram[33038] = 180;
// bram[33039] = 162;
// bram[33040] = 142;
// bram[33041] = 123;
// bram[33042] = 103;
// bram[33043] = 85;
// bram[33044] = 67;
// bram[33045] = 50;
// bram[33046] = 36;
// bram[33047] = 23;
// bram[33048] = 13;
// bram[33049] = 6;
// bram[33050] = 1;
// bram[33051] = 0;
// bram[33052] = 1;
// bram[33053] = 5;
// bram[33054] = 13;
// bram[33055] = 23;
// bram[33056] = 35;
// bram[33057] = 50;
// bram[33058] = 66;
// bram[33059] = 84;
// bram[33060] = 103;
// bram[33061] = 122;
// bram[33062] = 142;
// bram[33063] = 161;
// bram[33064] = 179;
// bram[33065] = 196;
// bram[33066] = 212;
// bram[33067] = 225;
// bram[33068] = 236;
// bram[33069] = 245;
// bram[33070] = 250;
// bram[33071] = 253;
// bram[33072] = 253;
// bram[33073] = 250;
// bram[33074] = 244;
// bram[33075] = 235;
// bram[33076] = 223;
// bram[33077] = 210;
// bram[33078] = 194;
// bram[33079] = 177;
// bram[33080] = 158;
// bram[33081] = 139;
// bram[33082] = 119;
// bram[33083] = 100;
// bram[33084] = 81;
// bram[33085] = 64;
// bram[33086] = 47;
// bram[33087] = 33;
// bram[33088] = 21;
// bram[33089] = 11;
// bram[33090] = 5;
// bram[33091] = 1;
// bram[33092] = 0;
// bram[33093] = 2;
// bram[33094] = 6;
// bram[33095] = 14;
// bram[33096] = 25;
// bram[33097] = 38;
// bram[33098] = 52;
// bram[33099] = 69;
// bram[33100] = 87;
// bram[33101] = 106;
// bram[33102] = 126;
// bram[33103] = 145;
// bram[33104] = 164;
// bram[33105] = 182;
// bram[33106] = 199;
// bram[33107] = 214;
// bram[33108] = 227;
// bram[33109] = 238;
// bram[33110] = 246;
// bram[33111] = 251;
// bram[33112] = 253;
// bram[33113] = 253;
// bram[33114] = 249;
// bram[33115] = 242;
// bram[33116] = 233;
// bram[33117] = 221;
// bram[33118] = 207;
// bram[33119] = 191;
// bram[33120] = 173;
// bram[33121] = 155;
// bram[33122] = 135;
// bram[33123] = 116;
// bram[33124] = 96;
// bram[33125] = 78;
// bram[33126] = 60;
// bram[33127] = 45;
// bram[33128] = 31;
// bram[33129] = 19;
// bram[33130] = 10;
// bram[33131] = 4;
// bram[33132] = 0;
// bram[33133] = 0;
// bram[33134] = 2;
// bram[33135] = 8;
// bram[33136] = 16;
// bram[33137] = 27;
// bram[33138] = 40;
// bram[33139] = 55;
// bram[33140] = 72;
// bram[33141] = 91;
// bram[33142] = 110;
// bram[33143] = 129;
// bram[33144] = 149;
// bram[33145] = 168;
// bram[33146] = 186;
// bram[33147] = 202;
// bram[33148] = 217;
// bram[33149] = 229;
// bram[33150] = 240;
// bram[33151] = 247;
// bram[33152] = 252;
// bram[33153] = 253;
// bram[33154] = 252;
// bram[33155] = 248;
// bram[33156] = 241;
// bram[33157] = 231;
// bram[33158] = 219;
// bram[33159] = 204;
// bram[33160] = 188;
// bram[33161] = 170;
// bram[33162] = 151;
// bram[33163] = 132;
// bram[33164] = 112;
// bram[33165] = 93;
// bram[33166] = 75;
// bram[33167] = 57;
// bram[33168] = 42;
// bram[33169] = 28;
// bram[33170] = 17;
// bram[33171] = 9;
// bram[33172] = 3;
// bram[33173] = 0;
// bram[33174] = 0;
// bram[33175] = 3;
// bram[33176] = 9;
// bram[33177] = 18;
// bram[33178] = 29;
// bram[33179] = 43;
// bram[33180] = 58;
// bram[33181] = 76;
// bram[33182] = 94;
// bram[33183] = 113;
// bram[33184] = 133;
// bram[33185] = 152;
// bram[33186] = 171;
// bram[33187] = 189;
// bram[33188] = 205;
// bram[33189] = 219;
// bram[33190] = 232;
// bram[33191] = 241;
// bram[33192] = 248;
// bram[33193] = 252;
// bram[33194] = 253;
// bram[33195] = 252;
// bram[33196] = 247;
// bram[33197] = 239;
// bram[33198] = 229;
// bram[33199] = 216;
// bram[33200] = 201;
// bram[33201] = 185;
// bram[33202] = 167;
// bram[33203] = 148;
// bram[33204] = 128;
// bram[33205] = 109;
// bram[33206] = 90;
// bram[33207] = 71;
// bram[33208] = 54;
// bram[33209] = 39;
// bram[33210] = 26;
// bram[33211] = 15;
// bram[33212] = 7;
// bram[33213] = 2;
// bram[33214] = 0;
// bram[33215] = 0;
// bram[33216] = 4;
// bram[33217] = 10;
// bram[33218] = 20;
// bram[33219] = 32;
// bram[33220] = 46;
// bram[33221] = 62;
// bram[33222] = 79;
// bram[33223] = 98;
// bram[33224] = 117;
// bram[33225] = 136;
// bram[33226] = 156;
// bram[33227] = 174;
// bram[33228] = 192;
// bram[33229] = 208;
// bram[33230] = 222;
// bram[33231] = 234;
// bram[33232] = 243;
// bram[33233] = 249;
// bram[33234] = 253;
// bram[33235] = 253;
// bram[33236] = 251;
// bram[33237] = 246;
// bram[33238] = 237;
// bram[33239] = 227;
// bram[33240] = 213;
// bram[33241] = 198;
// bram[33242] = 181;
// bram[33243] = 163;
// bram[33244] = 144;
// bram[33245] = 125;
// bram[33246] = 105;
// bram[33247] = 86;
// bram[33248] = 68;
// bram[33249] = 52;
// bram[33250] = 37;
// bram[33251] = 24;
// bram[33252] = 14;
// bram[33253] = 6;
// bram[33254] = 1;
// bram[33255] = 0;
// bram[33256] = 1;
// bram[33257] = 5;
// bram[33258] = 12;
// bram[33259] = 22;
// bram[33260] = 34;
// bram[33261] = 48;
// bram[33262] = 65;
// bram[33263] = 82;
// bram[33264] = 101;
// bram[33265] = 121;
// bram[33266] = 140;
// bram[33267] = 159;
// bram[33268] = 178;
// bram[33269] = 195;
// bram[33270] = 210;
// bram[33271] = 224;
// bram[33272] = 235;
// bram[33273] = 244;
// bram[33274] = 250;
// bram[33275] = 253;
// bram[33276] = 253;
// bram[33277] = 250;
// bram[33278] = 244;
// bram[33279] = 236;
// bram[33280] = 224;
// bram[33281] = 211;
// bram[33282] = 195;
// bram[33283] = 178;
// bram[33284] = 160;
// bram[33285] = 140;
// bram[33286] = 121;
// bram[33287] = 102;
// bram[33288] = 83;
// bram[33289] = 65;
// bram[33290] = 49;
// bram[33291] = 34;
// bram[33292] = 22;
// bram[33293] = 12;
// bram[33294] = 5;
// bram[33295] = 1;
// bram[33296] = 0;
// bram[33297] = 1;
// bram[33298] = 6;
// bram[33299] = 14;
// bram[33300] = 24;
// bram[33301] = 36;
// bram[33302] = 51;
// bram[33303] = 68;
// bram[33304] = 86;
// bram[33305] = 105;
// bram[33306] = 124;
// bram[33307] = 144;
// bram[33308] = 163;
// bram[33309] = 181;
// bram[33310] = 198;
// bram[33311] = 213;
// bram[33312] = 226;
// bram[33313] = 237;
// bram[33314] = 245;
// bram[33315] = 251;
// bram[33316] = 253;
// bram[33317] = 253;
// bram[33318] = 249;
// bram[33319] = 243;
// bram[33320] = 234;
// bram[33321] = 222;
// bram[33322] = 208;
// bram[33323] = 192;
// bram[33324] = 175;
// bram[33325] = 156;
// bram[33326] = 137;
// bram[33327] = 117;
// bram[33328] = 98;
// bram[33329] = 79;
// bram[33330] = 62;
// bram[33331] = 46;
// bram[33332] = 32;
// bram[33333] = 20;
// bram[33334] = 11;
// bram[33335] = 4;
// bram[33336] = 0;
// bram[33337] = 0;
// bram[33338] = 2;
// bram[33339] = 7;
// bram[33340] = 15;
// bram[33341] = 26;
// bram[33342] = 39;
// bram[33343] = 54;
// bram[33344] = 71;
// bram[33345] = 89;
// bram[33346] = 108;
// bram[33347] = 128;
// bram[33348] = 147;
// bram[33349] = 166;
// bram[33350] = 184;
// bram[33351] = 201;
// bram[33352] = 216;
// bram[33353] = 229;
// bram[33354] = 239;
// bram[33355] = 247;
// bram[33356] = 252;
// bram[33357] = 253;
// bram[33358] = 252;
// bram[33359] = 248;
// bram[33360] = 241;
// bram[33361] = 232;
// bram[33362] = 220;
// bram[33363] = 205;
// bram[33364] = 189;
// bram[33365] = 171;
// bram[33366] = 153;
// bram[33367] = 133;
// bram[33368] = 114;
// bram[33369] = 95;
// bram[33370] = 76;
// bram[33371] = 59;
// bram[33372] = 43;
// bram[33373] = 29;
// bram[33374] = 18;
// bram[33375] = 9;
// bram[33376] = 3;
// bram[33377] = 0;
// bram[33378] = 0;
// bram[33379] = 3;
// bram[33380] = 8;
// bram[33381] = 17;
// bram[33382] = 28;
// bram[33383] = 42;
// bram[33384] = 57;
// bram[33385] = 74;
// bram[33386] = 93;
// bram[33387] = 112;
// bram[33388] = 131;
// bram[33389] = 151;
// bram[33390] = 170;
// bram[33391] = 187;
// bram[33392] = 204;
// bram[33393] = 218;
// bram[33394] = 231;
// bram[33395] = 241;
// bram[33396] = 248;
// bram[33397] = 252;
// bram[33398] = 253;
// bram[33399] = 252;
// bram[33400] = 247;
// bram[33401] = 240;
// bram[33402] = 230;
// bram[33403] = 217;
// bram[33404] = 202;
// bram[33405] = 186;
// bram[33406] = 168;
// bram[33407] = 149;
// bram[33408] = 130;
// bram[33409] = 110;
// bram[33410] = 91;
// bram[33411] = 73;
// bram[33412] = 56;
// bram[33413] = 40;
// bram[33414] = 27;
// bram[33415] = 16;
// bram[33416] = 8;
// bram[33417] = 2;
// bram[33418] = 0;
// bram[33419] = 0;
// bram[33420] = 3;
// bram[33421] = 10;
// bram[33422] = 19;
// bram[33423] = 30;
// bram[33424] = 44;
// bram[33425] = 60;
// bram[33426] = 78;
// bram[33427] = 96;
// bram[33428] = 115;
// bram[33429] = 135;
// bram[33430] = 154;
// bram[33431] = 173;
// bram[33432] = 190;
// bram[33433] = 207;
// bram[33434] = 221;
// bram[33435] = 233;
// bram[33436] = 242;
// bram[33437] = 249;
// bram[33438] = 253;
// bram[33439] = 253;
// bram[33440] = 251;
// bram[33441] = 246;
// bram[33442] = 238;
// bram[33443] = 228;
// bram[33444] = 215;
// bram[33445] = 200;
// bram[33446] = 183;
// bram[33447] = 165;
// bram[33448] = 146;
// bram[33449] = 126;
// bram[33450] = 107;
// bram[33451] = 88;
// bram[33452] = 70;
// bram[33453] = 53;
// bram[33454] = 38;
// bram[33455] = 25;
// bram[33456] = 14;
// bram[33457] = 7;
// bram[33458] = 2;
// bram[33459] = 0;
// bram[33460] = 1;
// bram[33461] = 4;
// bram[33462] = 11;
// bram[33463] = 21;
// bram[33464] = 33;
// bram[33465] = 47;
// bram[33466] = 63;
// bram[33467] = 81;
// bram[33468] = 100;
// bram[33469] = 119;
// bram[33470] = 138;
// bram[33471] = 158;
// bram[33472] = 176;
// bram[33473] = 194;
// bram[33474] = 209;
// bram[33475] = 223;
// bram[33476] = 235;
// bram[33477] = 244;
// bram[33478] = 250;
// bram[33479] = 253;
// bram[33480] = 253;
// bram[33481] = 251;
// bram[33482] = 245;
// bram[33483] = 236;
// bram[33484] = 225;
// bram[33485] = 212;
// bram[33486] = 197;
// bram[33487] = 179;
// bram[33488] = 161;
// bram[33489] = 142;
// bram[33490] = 123;
// bram[33491] = 103;
// bram[33492] = 84;
// bram[33493] = 66;
// bram[33494] = 50;
// bram[33495] = 35;
// bram[33496] = 23;
// bram[33497] = 13;
// bram[33498] = 5;
// bram[33499] = 1;
// bram[33500] = 0;
// bram[33501] = 1;
// bram[33502] = 5;
// bram[33503] = 13;
// bram[33504] = 23;
// bram[33505] = 35;
// bram[33506] = 50;
// bram[33507] = 66;
// bram[33508] = 84;
// bram[33509] = 103;
// bram[33510] = 123;
// bram[33511] = 142;
// bram[33512] = 161;
// bram[33513] = 179;
// bram[33514] = 197;
// bram[33515] = 212;
// bram[33516] = 225;
// bram[33517] = 236;
// bram[33518] = 245;
// bram[33519] = 251;
// bram[33520] = 253;
// bram[33521] = 253;
// bram[33522] = 250;
// bram[33523] = 244;
// bram[33524] = 235;
// bram[33525] = 223;
// bram[33526] = 209;
// bram[33527] = 194;
// bram[33528] = 176;
// bram[33529] = 158;
// bram[33530] = 138;
// bram[33531] = 119;
// bram[33532] = 100;
// bram[33533] = 81;
// bram[33534] = 63;
// bram[33535] = 47;
// bram[33536] = 33;
// bram[33537] = 21;
// bram[33538] = 11;
// bram[33539] = 4;
// bram[33540] = 1;
// bram[33541] = 0;
// bram[33542] = 2;
// bram[33543] = 7;
// bram[33544] = 14;
// bram[33545] = 25;
// bram[33546] = 38;
// bram[33547] = 53;
// bram[33548] = 70;
// bram[33549] = 88;
// bram[33550] = 107;
// bram[33551] = 126;
// bram[33552] = 146;
// bram[33553] = 165;
// bram[33554] = 183;
// bram[33555] = 200;
// bram[33556] = 215;
// bram[33557] = 228;
// bram[33558] = 238;
// bram[33559] = 246;
// bram[33560] = 251;
// bram[33561] = 253;
// bram[33562] = 253;
// bram[33563] = 249;
// bram[33564] = 242;
// bram[33565] = 233;
// bram[33566] = 221;
// bram[33567] = 207;
// bram[33568] = 190;
// bram[33569] = 173;
// bram[33570] = 154;
// bram[33571] = 135;
// bram[33572] = 115;
// bram[33573] = 96;
// bram[33574] = 78;
// bram[33575] = 60;
// bram[33576] = 44;
// bram[33577] = 30;
// bram[33578] = 19;
// bram[33579] = 10;
// bram[33580] = 3;
// bram[33581] = 0;
// bram[33582] = 0;
// bram[33583] = 2;
// bram[33584] = 8;
// bram[33585] = 16;
// bram[33586] = 27;
// bram[33587] = 40;
// bram[33588] = 56;
// bram[33589] = 73;
// bram[33590] = 91;
// bram[33591] = 110;
// bram[33592] = 130;
// bram[33593] = 149;
// bram[33594] = 168;
// bram[33595] = 186;
// bram[33596] = 202;
// bram[33597] = 217;
// bram[33598] = 230;
// bram[33599] = 240;
// bram[33600] = 247;
// bram[33601] = 252;
// bram[33602] = 253;
// bram[33603] = 252;
// bram[33604] = 248;
// bram[33605] = 241;
// bram[33606] = 231;
// bram[33607] = 218;
// bram[33608] = 204;
// bram[33609] = 187;
// bram[33610] = 170;
// bram[33611] = 151;
// bram[33612] = 131;
// bram[33613] = 112;
// bram[33614] = 93;
// bram[33615] = 74;
// bram[33616] = 57;
// bram[33617] = 42;
// bram[33618] = 28;
// bram[33619] = 17;
// bram[33620] = 8;
// bram[33621] = 3;
// bram[33622] = 0;
// bram[33623] = 0;
// bram[33624] = 3;
// bram[33625] = 9;
// bram[33626] = 18;
// bram[33627] = 29;
// bram[33628] = 43;
// bram[33629] = 59;
// bram[33630] = 76;
// bram[33631] = 95;
// bram[33632] = 114;
// bram[33633] = 133;
// bram[33634] = 153;
// bram[33635] = 171;
// bram[33636] = 189;
// bram[33637] = 205;
// bram[33638] = 220;
// bram[33639] = 232;
// bram[33640] = 241;
// bram[33641] = 248;
// bram[33642] = 252;
// bram[33643] = 253;
// bram[33644] = 252;
// bram[33645] = 247;
// bram[33646] = 239;
// bram[33647] = 229;
// bram[33648] = 216;
// bram[33649] = 201;
// bram[33650] = 184;
// bram[33651] = 166;
// bram[33652] = 147;
// bram[33653] = 128;
// bram[33654] = 108;
// bram[33655] = 89;
// bram[33656] = 71;
// bram[33657] = 54;
// bram[33658] = 39;
// bram[33659] = 26;
// bram[33660] = 15;
// bram[33661] = 7;
// bram[33662] = 2;
// bram[33663] = 0;
// bram[33664] = 0;
// bram[33665] = 4;
// bram[33666] = 11;
// bram[33667] = 20;
// bram[33668] = 32;
// bram[33669] = 46;
// bram[33670] = 62;
// bram[33671] = 79;
// bram[33672] = 98;
// bram[33673] = 117;
// bram[33674] = 137;
// bram[33675] = 156;
// bram[33676] = 175;
// bram[33677] = 192;
// bram[33678] = 208;
// bram[33679] = 222;
// bram[33680] = 234;
// bram[33681] = 243;
// bram[33682] = 249;
// bram[33683] = 253;
// bram[33684] = 253;
// bram[33685] = 251;
// bram[33686] = 245;
// bram[33687] = 237;
// bram[33688] = 226;
// bram[33689] = 213;
// bram[33690] = 198;
// bram[33691] = 181;
// bram[33692] = 163;
// bram[33693] = 144;
// bram[33694] = 124;
// bram[33695] = 105;
// bram[33696] = 86;
// bram[33697] = 68;
// bram[33698] = 51;
// bram[33699] = 36;
// bram[33700] = 24;
// bram[33701] = 14;
// bram[33702] = 6;
// bram[33703] = 1;
// bram[33704] = 0;
// bram[33705] = 1;
// bram[33706] = 5;
// bram[33707] = 12;
// bram[33708] = 22;
// bram[33709] = 34;
// bram[33710] = 49;
// bram[33711] = 65;
// bram[33712] = 83;
// bram[33713] = 102;
// bram[33714] = 121;
// bram[33715] = 140;
// bram[33716] = 160;
// bram[33717] = 178;
// bram[33718] = 195;
// bram[33719] = 211;
// bram[33720] = 224;
// bram[33721] = 236;
// bram[33722] = 244;
// bram[33723] = 250;
// bram[33724] = 253;
// bram[33725] = 253;
// bram[33726] = 250;
// bram[33727] = 244;
// bram[33728] = 235;
// bram[33729] = 224;
// bram[33730] = 210;
// bram[33731] = 195;
// bram[33732] = 178;
// bram[33733] = 159;
// bram[33734] = 140;
// bram[33735] = 121;
// bram[33736] = 101;
// bram[33737] = 82;
// bram[33738] = 65;
// bram[33739] = 48;
// bram[33740] = 34;
// bram[33741] = 22;
// bram[33742] = 12;
// bram[33743] = 5;
// bram[33744] = 1;
// bram[33745] = 0;
// bram[33746] = 1;
// bram[33747] = 6;
// bram[33748] = 14;
// bram[33749] = 24;
// bram[33750] = 37;
// bram[33751] = 52;
// bram[33752] = 68;
// bram[33753] = 86;
// bram[33754] = 105;
// bram[33755] = 125;
// bram[33756] = 144;
// bram[33757] = 163;
// bram[33758] = 181;
// bram[33759] = 198;
// bram[33760] = 213;
// bram[33761] = 227;
// bram[33762] = 237;
// bram[33763] = 246;
// bram[33764] = 251;
// bram[33765] = 253;
// bram[33766] = 253;
// bram[33767] = 249;
// bram[33768] = 243;
// bram[33769] = 234;
// bram[33770] = 222;
// bram[33771] = 208;
// bram[33772] = 192;
// bram[33773] = 174;
// bram[33774] = 156;
// bram[33775] = 136;
// bram[33776] = 117;
// bram[33777] = 98;
// bram[33778] = 79;
// bram[33779] = 62;
// bram[33780] = 46;
// bram[33781] = 32;
// bram[33782] = 20;
// bram[33783] = 10;
// bram[33784] = 4;
// bram[33785] = 0;
// bram[33786] = 0;
// bram[33787] = 2;
// bram[33788] = 7;
// bram[33789] = 15;
// bram[33790] = 26;
// bram[33791] = 39;
// bram[33792] = 54;
// bram[33793] = 71;
// bram[33794] = 90;
// bram[33795] = 109;
// bram[33796] = 128;
// bram[33797] = 148;
// bram[33798] = 167;
// bram[33799] = 185;
// bram[33800] = 201;
// bram[33801] = 216;
// bram[33802] = 229;
// bram[33803] = 239;
// bram[33804] = 247;
// bram[33805] = 252;
// bram[33806] = 253;
// bram[33807] = 252;
// bram[33808] = 248;
// bram[33809] = 241;
// bram[33810] = 232;
// bram[33811] = 219;
// bram[33812] = 205;
// bram[33813] = 189;
// bram[33814] = 171;
// bram[33815] = 152;
// bram[33816] = 133;
// bram[33817] = 113;
// bram[33818] = 94;
// bram[33819] = 76;
// bram[33820] = 58;
// bram[33821] = 43;
// bram[33822] = 29;
// bram[33823] = 18;
// bram[33824] = 9;
// bram[33825] = 3;
// bram[33826] = 0;
// bram[33827] = 0;
// bram[33828] = 3;
// bram[33829] = 9;
// bram[33830] = 17;
// bram[33831] = 28;
// bram[33832] = 42;
// bram[33833] = 57;
// bram[33834] = 75;
// bram[33835] = 93;
// bram[33836] = 112;
// bram[33837] = 132;
// bram[33838] = 151;
// bram[33839] = 170;
// bram[33840] = 188;
// bram[33841] = 204;
// bram[33842] = 219;
// bram[33843] = 231;
// bram[33844] = 241;
// bram[33845] = 248;
// bram[33846] = 252;
// bram[33847] = 253;
// bram[33848] = 252;
// bram[33849] = 247;
// bram[33850] = 240;
// bram[33851] = 229;
// bram[33852] = 217;
// bram[33853] = 202;
// bram[33854] = 186;
// bram[33855] = 168;
// bram[33856] = 149;
// bram[33857] = 129;
// bram[33858] = 110;
// bram[33859] = 91;
// bram[33860] = 72;
// bram[33861] = 55;
// bram[33862] = 40;
// bram[33863] = 27;
// bram[33864] = 16;
// bram[33865] = 8;
// bram[33866] = 2;
// bram[33867] = 0;
// bram[33868] = 0;
// bram[33869] = 4;
// bram[33870] = 10;
// bram[33871] = 19;
// bram[33872] = 31;
// bram[33873] = 45;
// bram[33874] = 60;
// bram[33875] = 78;
// bram[33876] = 96;
// bram[33877] = 116;
// bram[33878] = 135;
// bram[33879] = 155;
// bram[33880] = 173;
// bram[33881] = 191;
// bram[33882] = 207;
// bram[33883] = 221;
// bram[33884] = 233;
// bram[33885] = 242;
// bram[33886] = 249;
// bram[33887] = 253;
// bram[33888] = 253;
// bram[33889] = 251;
// bram[33890] = 246;
// bram[33891] = 238;
// bram[33892] = 227;
// bram[33893] = 214;
// bram[33894] = 199;
// bram[33895] = 182;
// bram[33896] = 164;
// bram[33897] = 145;
// bram[33898] = 126;
// bram[33899] = 106;
// bram[33900] = 87;
// bram[33901] = 69;
// bram[33902] = 52;
// bram[33903] = 38;
// bram[33904] = 25;
// bram[33905] = 14;
// bram[33906] = 6;
// bram[33907] = 2;
// bram[33908] = 0;
// bram[33909] = 1;
// bram[33910] = 5;
// bram[33911] = 11;
// bram[33912] = 21;
// bram[33913] = 33;
// bram[33914] = 47;
// bram[33915] = 64;
// bram[33916] = 81;
// bram[33917] = 100;
// bram[33918] = 119;
// bram[33919] = 139;
// bram[33920] = 158;
// bram[33921] = 177;
// bram[33922] = 194;
// bram[33923] = 210;
// bram[33924] = 223;
// bram[33925] = 235;
// bram[33926] = 244;
// bram[33927] = 250;
// bram[33928] = 253;
// bram[33929] = 253;
// bram[33930] = 250;
// bram[33931] = 245;
// bram[33932] = 236;
// bram[33933] = 225;
// bram[33934] = 212;
// bram[33935] = 196;
// bram[33936] = 179;
// bram[33937] = 161;
// bram[33938] = 142;
// bram[33939] = 122;
// bram[33940] = 103;
// bram[33941] = 84;
// bram[33942] = 66;
// bram[33943] = 50;
// bram[33944] = 35;
// bram[33945] = 23;
// bram[33946] = 13;
// bram[33947] = 5;
// bram[33948] = 1;
// bram[33949] = 0;
// bram[33950] = 1;
// bram[33951] = 6;
// bram[33952] = 13;
// bram[33953] = 23;
// bram[33954] = 36;
// bram[33955] = 50;
// bram[33956] = 67;
// bram[33957] = 85;
// bram[33958] = 103;
// bram[33959] = 123;
// bram[33960] = 142;
// bram[33961] = 162;
// bram[33962] = 180;
// bram[33963] = 197;
// bram[33964] = 212;
// bram[33965] = 226;
// bram[33966] = 237;
// bram[33967] = 245;
// bram[33968] = 251;
// bram[33969] = 253;
// bram[33970] = 253;
// bram[33971] = 250;
// bram[33972] = 243;
// bram[33973] = 234;
// bram[33974] = 223;
// bram[33975] = 209;
// bram[33976] = 193;
// bram[33977] = 176;
// bram[33978] = 157;
// bram[33979] = 138;
// bram[33980] = 119;
// bram[33981] = 99;
// bram[33982] = 80;
// bram[33983] = 63;
// bram[33984] = 47;
// bram[33985] = 33;
// bram[33986] = 21;
// bram[33987] = 11;
// bram[33988] = 4;
// bram[33989] = 0;
// bram[33990] = 0;
// bram[33991] = 2;
// bram[33992] = 7;
// bram[33993] = 15;
// bram[33994] = 25;
// bram[33995] = 38;
// bram[33996] = 53;
// bram[33997] = 70;
// bram[33998] = 88;
// bram[33999] = 107;
// bram[34000] = 126;
// bram[34001] = 146;
// bram[34002] = 165;
// bram[34003] = 183;
// bram[34004] = 200;
// bram[34005] = 215;
// bram[34006] = 228;
// bram[34007] = 238;
// bram[34008] = 246;
// bram[34009] = 251;
// bram[34010] = 253;
// bram[34011] = 253;
// bram[34012] = 249;
// bram[34013] = 242;
// bram[34014] = 232;
// bram[34015] = 220;
// bram[34016] = 206;
// bram[34017] = 190;
// bram[34018] = 173;
// bram[34019] = 154;
// bram[34020] = 134;
// bram[34021] = 115;
// bram[34022] = 96;
// bram[34023] = 77;
// bram[34024] = 60;
// bram[34025] = 44;
// bram[34026] = 30;
// bram[34027] = 19;
// bram[34028] = 10;
// bram[34029] = 3;
// bram[34030] = 0;
// bram[34031] = 0;
// bram[34032] = 2;
// bram[34033] = 8;
// bram[34034] = 16;
// bram[34035] = 27;
// bram[34036] = 41;
// bram[34037] = 56;
// bram[34038] = 73;
// bram[34039] = 91;
// bram[34040] = 111;
// bram[34041] = 130;
// bram[34042] = 150;
// bram[34043] = 168;
// bram[34044] = 186;
// bram[34045] = 203;
// bram[34046] = 217;
// bram[34047] = 230;
// bram[34048] = 240;
// bram[34049] = 247;
// bram[34050] = 252;
// bram[34051] = 253;
// bram[34052] = 252;
// bram[34053] = 248;
// bram[34054] = 240;
// bram[34055] = 230;
// bram[34056] = 218;
// bram[34057] = 203;
// bram[34058] = 187;
// bram[34059] = 169;
// bram[34060] = 150;
// bram[34061] = 131;
// bram[34062] = 111;
// bram[34063] = 92;
// bram[34064] = 74;
// bram[34065] = 57;
// bram[34066] = 41;
// bram[34067] = 28;
// bram[34068] = 17;
// bram[34069] = 8;
// bram[34070] = 3;
// bram[34071] = 0;
// bram[34072] = 0;
// bram[34073] = 3;
// bram[34074] = 9;
// bram[34075] = 18;
// bram[34076] = 30;
// bram[34077] = 43;
// bram[34078] = 59;
// bram[34079] = 76;
// bram[34080] = 95;
// bram[34081] = 114;
// bram[34082] = 134;
// bram[34083] = 153;
// bram[34084] = 172;
// bram[34085] = 189;
// bram[34086] = 206;
// bram[34087] = 220;
// bram[34088] = 232;
// bram[34089] = 242;
// bram[34090] = 248;
// bram[34091] = 252;
// bram[34092] = 253;
// bram[34093] = 251;
// bram[34094] = 247;
// bram[34095] = 239;
// bram[34096] = 228;
// bram[34097] = 215;
// bram[34098] = 201;
// bram[34099] = 184;
// bram[34100] = 166;
// bram[34101] = 147;
// bram[34102] = 127;
// bram[34103] = 108;
// bram[34104] = 89;
// bram[34105] = 71;
// bram[34106] = 54;
// bram[34107] = 39;
// bram[34108] = 26;
// bram[34109] = 15;
// bram[34110] = 7;
// bram[34111] = 2;
// bram[34112] = 0;
// bram[34113] = 0;
// bram[34114] = 4;
// bram[34115] = 11;
// bram[34116] = 20;
// bram[34117] = 32;
// bram[34118] = 46;
// bram[34119] = 62;
// bram[34120] = 80;
// bram[34121] = 98;
// bram[34122] = 118;
// bram[34123] = 137;
// bram[34124] = 157;
// bram[34125] = 175;
// bram[34126] = 193;
// bram[34127] = 208;
// bram[34128] = 222;
// bram[34129] = 234;
// bram[34130] = 243;
// bram[34131] = 249;
// bram[34132] = 253;
// bram[34133] = 253;
// bram[34134] = 251;
// bram[34135] = 245;
// bram[34136] = 237;
// bram[34137] = 226;
// bram[34138] = 213;
// bram[34139] = 198;
// bram[34140] = 181;
// bram[34141] = 162;
// bram[34142] = 143;
// bram[34143] = 124;
// bram[34144] = 104;
// bram[34145] = 85;
// bram[34146] = 67;
// bram[34147] = 51;
// bram[34148] = 36;
// bram[34149] = 24;
// bram[34150] = 13;
// bram[34151] = 6;
// bram[34152] = 1;
// bram[34153] = 0;
// bram[34154] = 1;
// bram[34155] = 5;
// bram[34156] = 12;
// bram[34157] = 22;
// bram[34158] = 34;
// bram[34159] = 49;
// bram[34160] = 65;
// bram[34161] = 83;
// bram[34162] = 102;
// bram[34163] = 121;
// bram[34164] = 141;
// bram[34165] = 160;
// bram[34166] = 178;
// bram[34167] = 196;
// bram[34168] = 211;
// bram[34169] = 225;
// bram[34170] = 236;
// bram[34171] = 244;
// bram[34172] = 250;
// bram[34173] = 253;
// bram[34174] = 253;
// bram[34175] = 250;
// bram[34176] = 244;
// bram[34177] = 235;
// bram[34178] = 224;
// bram[34179] = 210;
// bram[34180] = 195;
// bram[34181] = 177;
// bram[34182] = 159;
// bram[34183] = 140;
// bram[34184] = 120;
// bram[34185] = 101;
// bram[34186] = 82;
// bram[34187] = 64;
// bram[34188] = 48;
// bram[34189] = 34;
// bram[34190] = 21;
// bram[34191] = 12;
// bram[34192] = 5;
// bram[34193] = 1;
// bram[34194] = 0;
// bram[34195] = 1;
// bram[34196] = 6;
// bram[34197] = 14;
// bram[34198] = 24;
// bram[34199] = 37;
// bram[34200] = 52;
// bram[34201] = 68;
// bram[34202] = 86;
// bram[34203] = 105;
// bram[34204] = 125;
// bram[34205] = 144;
// bram[34206] = 163;
// bram[34207] = 182;
// bram[34208] = 199;
// bram[34209] = 214;
// bram[34210] = 227;
// bram[34211] = 238;
// bram[34212] = 246;
// bram[34213] = 251;
// bram[34214] = 253;
// bram[34215] = 253;
// bram[34216] = 249;
// bram[34217] = 243;
// bram[34218] = 233;
// bram[34219] = 221;
// bram[34220] = 207;
// bram[34221] = 191;
// bram[34222] = 174;
// bram[34223] = 155;
// bram[34224] = 136;
// bram[34225] = 117;
// bram[34226] = 97;
// bram[34227] = 79;
// bram[34228] = 61;
// bram[34229] = 45;
// bram[34230] = 31;
// bram[34231] = 19;
// bram[34232] = 10;
// bram[34233] = 4;
// bram[34234] = 0;
// bram[34235] = 0;
// bram[34236] = 2;
// bram[34237] = 7;
// bram[34238] = 16;
// bram[34239] = 26;
// bram[34240] = 40;
// bram[34241] = 55;
// bram[34242] = 72;
// bram[34243] = 90;
// bram[34244] = 109;
// bram[34245] = 128;
// bram[34246] = 148;
// bram[34247] = 167;
// bram[34248] = 185;
// bram[34249] = 201;
// bram[34250] = 216;
// bram[34251] = 229;
// bram[34252] = 239;
// bram[34253] = 247;
// bram[34254] = 252;
// bram[34255] = 253;
// bram[34256] = 252;
// bram[34257] = 248;
// bram[34258] = 241;
// bram[34259] = 231;
// bram[34260] = 219;
// bram[34261] = 205;
// bram[34262] = 188;
// bram[34263] = 171;
// bram[34264] = 152;
// bram[34265] = 132;
// bram[34266] = 113;
// bram[34267] = 94;
// bram[34268] = 75;
// bram[34269] = 58;
// bram[34270] = 43;
// bram[34271] = 29;
// bram[34272] = 18;
// bram[34273] = 9;
// bram[34274] = 3;
// bram[34275] = 0;
// bram[34276] = 0;
// bram[34277] = 3;
// bram[34278] = 9;
// bram[34279] = 17;
// bram[34280] = 29;
// bram[34281] = 42;
// bram[34282] = 58;
// bram[34283] = 75;
// bram[34284] = 93;
// bram[34285] = 113;
// bram[34286] = 132;
// bram[34287] = 151;
// bram[34288] = 170;
// bram[34289] = 188;
// bram[34290] = 204;
// bram[34291] = 219;
// bram[34292] = 231;
// bram[34293] = 241;
// bram[34294] = 248;
// bram[34295] = 252;
// bram[34296] = 253;
// bram[34297] = 252;
// bram[34298] = 247;
// bram[34299] = 239;
// bram[34300] = 229;
// bram[34301] = 217;
// bram[34302] = 202;
// bram[34303] = 185;
// bram[34304] = 167;
// bram[34305] = 148;
// bram[34306] = 129;
// bram[34307] = 109;
// bram[34308] = 90;
// bram[34309] = 72;
// bram[34310] = 55;
// bram[34311] = 40;
// bram[34312] = 27;
// bram[34313] = 16;
// bram[34314] = 8;
// bram[34315] = 2;
// bram[34316] = 0;
// bram[34317] = 0;
// bram[34318] = 4;
// bram[34319] = 10;
// bram[34320] = 19;
// bram[34321] = 31;
// bram[34322] = 45;
// bram[34323] = 61;
// bram[34324] = 78;
// bram[34325] = 97;
// bram[34326] = 116;
// bram[34327] = 136;
// bram[34328] = 155;
// bram[34329] = 174;
// bram[34330] = 191;
// bram[34331] = 207;
// bram[34332] = 221;
// bram[34333] = 233;
// bram[34334] = 242;
// bram[34335] = 249;
// bram[34336] = 253;
// bram[34337] = 253;
// bram[34338] = 251;
// bram[34339] = 246;
// bram[34340] = 238;
// bram[34341] = 227;
// bram[34342] = 214;
// bram[34343] = 199;
// bram[34344] = 182;
// bram[34345] = 164;
// bram[34346] = 145;
// bram[34347] = 125;
// bram[34348] = 106;
// bram[34349] = 87;
// bram[34350] = 69;
// bram[34351] = 52;
// bram[34352] = 37;
// bram[34353] = 24;
// bram[34354] = 14;
// bram[34355] = 6;
// bram[34356] = 1;
// bram[34357] = 0;
// bram[34358] = 1;
// bram[34359] = 5;
// bram[34360] = 12;
// bram[34361] = 21;
// bram[34362] = 33;
// bram[34363] = 48;
// bram[34364] = 64;
// bram[34365] = 82;
// bram[34366] = 100;
// bram[34367] = 120;
// bram[34368] = 139;
// bram[34369] = 158;
// bram[34370] = 177;
// bram[34371] = 194;
// bram[34372] = 210;
// bram[34373] = 224;
// bram[34374] = 235;
// bram[34375] = 244;
// bram[34376] = 250;
// bram[34377] = 253;
// bram[34378] = 253;
// bram[34379] = 250;
// bram[34380] = 245;
// bram[34381] = 236;
// bram[34382] = 225;
// bram[34383] = 211;
// bram[34384] = 196;
// bram[34385] = 179;
// bram[34386] = 160;
// bram[34387] = 141;
// bram[34388] = 122;
// bram[34389] = 102;
// bram[34390] = 83;
// bram[34391] = 66;
// bram[34392] = 49;
// bram[34393] = 35;
// bram[34394] = 22;
// bram[34395] = 12;
// bram[34396] = 5;
// bram[34397] = 1;
// bram[34398] = 0;
// bram[34399] = 1;
// bram[34400] = 6;
// bram[34401] = 13;
// bram[34402] = 23;
// bram[34403] = 36;
// bram[34404] = 51;
// bram[34405] = 67;
// bram[34406] = 85;
// bram[34407] = 104;
// bram[34408] = 123;
// bram[34409] = 143;
// bram[34410] = 162;
// bram[34411] = 180;
// bram[34412] = 197;
// bram[34413] = 213;
// bram[34414] = 226;
// bram[34415] = 237;
// bram[34416] = 245;
// bram[34417] = 251;
// bram[34418] = 253;
// bram[34419] = 253;
// bram[34420] = 250;
// bram[34421] = 243;
// bram[34422] = 234;
// bram[34423] = 223;
// bram[34424] = 209;
// bram[34425] = 193;
// bram[34426] = 175;
// bram[34427] = 157;
// bram[34428] = 138;
// bram[34429] = 118;
// bram[34430] = 99;
// bram[34431] = 80;
// bram[34432] = 63;
// bram[34433] = 46;
// bram[34434] = 32;
// bram[34435] = 20;
// bram[34436] = 11;
// bram[34437] = 4;
// bram[34438] = 0;
// bram[34439] = 0;
// bram[34440] = 2;
// bram[34441] = 7;
// bram[34442] = 15;
// bram[34443] = 25;
// bram[34444] = 38;
// bram[34445] = 53;
// bram[34446] = 70;
// bram[34447] = 88;
// bram[34448] = 107;
// bram[34449] = 127;
// bram[34450] = 146;
// bram[34451] = 165;
// bram[34452] = 183;
// bram[34453] = 200;
// bram[34454] = 215;
// bram[34455] = 228;
// bram[34456] = 239;
// bram[34457] = 246;
// bram[34458] = 251;
// bram[34459] = 253;
// bram[34460] = 252;
// bram[34461] = 249;
// bram[34462] = 242;
// bram[34463] = 232;
// bram[34464] = 220;
// bram[34465] = 206;
// bram[34466] = 190;
// bram[34467] = 172;
// bram[34468] = 153;
// bram[34469] = 134;
// bram[34470] = 115;
// bram[34471] = 95;
// bram[34472] = 77;
// bram[34473] = 59;
// bram[34474] = 44;
// bram[34475] = 30;
// bram[34476] = 18;
// bram[34477] = 9;
// bram[34478] = 3;
// bram[34479] = 0;
// bram[34480] = 0;
// bram[34481] = 2;
// bram[34482] = 8;
// bram[34483] = 17;
// bram[34484] = 28;
// bram[34485] = 41;
// bram[34486] = 56;
// bram[34487] = 74;
// bram[34488] = 92;
// bram[34489] = 111;
// bram[34490] = 130;
// bram[34491] = 150;
// bram[34492] = 169;
// bram[34493] = 187;
// bram[34494] = 203;
// bram[34495] = 218;
// bram[34496] = 230;
// bram[34497] = 240;
// bram[34498] = 248;
// bram[34499] = 252;
// bram[34500] = 254;
// bram[34501] = 252;
// bram[34502] = 248;
// bram[34503] = 240;
// bram[34504] = 230;
// bram[34505] = 218;
// bram[34506] = 203;
// bram[34507] = 187;
// bram[34508] = 169;
// bram[34509] = 150;
// bram[34510] = 130;
// bram[34511] = 111;
// bram[34512] = 92;
// bram[34513] = 74;
// bram[34514] = 56;
// bram[34515] = 41;
// bram[34516] = 28;
// bram[34517] = 17;
// bram[34518] = 8;
// bram[34519] = 2;
// bram[34520] = 0;
// bram[34521] = 0;
// bram[34522] = 3;
// bram[34523] = 9;
// bram[34524] = 18;
// bram[34525] = 30;
// bram[34526] = 44;
// bram[34527] = 59;
// bram[34528] = 77;
// bram[34529] = 95;
// bram[34530] = 115;
// bram[34531] = 134;
// bram[34532] = 153;
// bram[34533] = 172;
// bram[34534] = 190;
// bram[34535] = 206;
// bram[34536] = 220;
// bram[34537] = 232;
// bram[34538] = 242;
// bram[34539] = 249;
// bram[34540] = 252;
// bram[34541] = 253;
// bram[34542] = 251;
// bram[34543] = 246;
// bram[34544] = 239;
// bram[34545] = 228;
// bram[34546] = 215;
// bram[34547] = 200;
// bram[34548] = 183;
// bram[34549] = 165;
// bram[34550] = 146;
// bram[34551] = 127;
// bram[34552] = 107;
// bram[34553] = 88;
// bram[34554] = 70;
// bram[34555] = 53;
// bram[34556] = 38;
// bram[34557] = 25;
// bram[34558] = 15;
// bram[34559] = 7;
// bram[34560] = 2;
// bram[34561] = 0;
// bram[34562] = 0;
// bram[34563] = 4;
// bram[34564] = 11;
// bram[34565] = 20;
// bram[34566] = 32;
// bram[34567] = 46;
// bram[34568] = 63;
// bram[34569] = 80;
// bram[34570] = 99;
// bram[34571] = 118;
// bram[34572] = 138;
// bram[34573] = 157;
// bram[34574] = 175;
// bram[34575] = 193;
// bram[34576] = 209;
// bram[34577] = 223;
// bram[34578] = 234;
// bram[34579] = 243;
// bram[34580] = 250;
// bram[34581] = 253;
// bram[34582] = 253;
// bram[34583] = 251;
// bram[34584] = 245;
// bram[34585] = 237;
// bram[34586] = 226;
// bram[34587] = 213;
// bram[34588] = 197;
// bram[34589] = 180;
// bram[34590] = 162;
// bram[34591] = 143;
// bram[34592] = 123;
// bram[34593] = 104;
// bram[34594] = 85;
// bram[34595] = 67;
// bram[34596] = 51;
// bram[34597] = 36;
// bram[34598] = 23;
// bram[34599] = 13;
// bram[34600] = 6;
// bram[34601] = 1;
// bram[34602] = 0;
// bram[34603] = 1;
// bram[34604] = 5;
// bram[34605] = 12;
// bram[34606] = 22;
// bram[34607] = 35;
// bram[34608] = 49;
// bram[34609] = 66;
// bram[34610] = 83;
// bram[34611] = 102;
// bram[34612] = 122;
// bram[34613] = 141;
// bram[34614] = 160;
// bram[34615] = 179;
// bram[34616] = 196;
// bram[34617] = 211;
// bram[34618] = 225;
// bram[34619] = 236;
// bram[34620] = 245;
// bram[34621] = 250;
// bram[34622] = 253;
// bram[34623] = 253;
// bram[34624] = 250;
// bram[34625] = 244;
// bram[34626] = 235;
// bram[34627] = 224;
// bram[34628] = 210;
// bram[34629] = 194;
// bram[34630] = 177;
// bram[34631] = 158;
// bram[34632] = 139;
// bram[34633] = 120;
// bram[34634] = 100;
// bram[34635] = 82;
// bram[34636] = 64;
// bram[34637] = 48;
// bram[34638] = 33;
// bram[34639] = 21;
// bram[34640] = 12;
// bram[34641] = 5;
// bram[34642] = 1;
// bram[34643] = 0;
// bram[34644] = 1;
// bram[34645] = 6;
// bram[34646] = 14;
// bram[34647] = 24;
// bram[34648] = 37;
// bram[34649] = 52;
// bram[34650] = 69;
// bram[34651] = 87;
// bram[34652] = 106;
// bram[34653] = 125;
// bram[34654] = 145;
// bram[34655] = 164;
// bram[34656] = 182;
// bram[34657] = 199;
// bram[34658] = 214;
// bram[34659] = 227;
// bram[34660] = 238;
// bram[34661] = 246;
// bram[34662] = 251;
// bram[34663] = 253;
// bram[34664] = 253;
// bram[34665] = 249;
// bram[34666] = 242;
// bram[34667] = 233;
// bram[34668] = 221;
// bram[34669] = 207;
// bram[34670] = 191;
// bram[34671] = 174;
// bram[34672] = 155;
// bram[34673] = 136;
// bram[34674] = 116;
// bram[34675] = 97;
// bram[34676] = 78;
// bram[34677] = 61;
// bram[34678] = 45;
// bram[34679] = 31;
// bram[34680] = 19;
// bram[34681] = 10;
// bram[34682] = 4;
// bram[34683] = 0;
// bram[34684] = 0;
// bram[34685] = 2;
// bram[34686] = 8;
// bram[34687] = 16;
// bram[34688] = 27;
// bram[34689] = 40;
// bram[34690] = 55;
// bram[34691] = 72;
// bram[34692] = 90;
// bram[34693] = 109;
// bram[34694] = 129;
// bram[34695] = 148;
// bram[34696] = 167;
// bram[34697] = 185;
// bram[34698] = 202;
// bram[34699] = 217;
// bram[34700] = 229;
// bram[34701] = 239;
// bram[34702] = 247;
// bram[34703] = 252;
// bram[34704] = 253;
// bram[34705] = 252;
// bram[34706] = 248;
// bram[34707] = 241;
// bram[34708] = 231;
// bram[34709] = 219;
// bram[34710] = 204;
// bram[34711] = 188;
// bram[34712] = 170;
// bram[34713] = 151;
// bram[34714] = 132;
// bram[34715] = 113;
// bram[34716] = 93;
// bram[34717] = 75;
// bram[34718] = 58;
// bram[34719] = 42;
// bram[34720] = 29;
// bram[34721] = 17;
// bram[34722] = 9;
// bram[34723] = 3;
// bram[34724] = 0;
// bram[34725] = 0;
// bram[34726] = 3;
// bram[34727] = 9;
// bram[34728] = 18;
// bram[34729] = 29;
// bram[34730] = 43;
// bram[34731] = 58;
// bram[34732] = 75;
// bram[34733] = 94;
// bram[34734] = 113;
// bram[34735] = 132;
// bram[34736] = 152;
// bram[34737] = 171;
// bram[34738] = 188;
// bram[34739] = 205;
// bram[34740] = 219;
// bram[34741] = 231;
// bram[34742] = 241;
// bram[34743] = 248;
// bram[34744] = 252;
// bram[34745] = 253;
// bram[34746] = 252;
// bram[34747] = 247;
// bram[34748] = 239;
// bram[34749] = 229;
// bram[34750] = 216;
// bram[34751] = 201;
// bram[34752] = 185;
// bram[34753] = 167;
// bram[34754] = 148;
// bram[34755] = 128;
// bram[34756] = 109;
// bram[34757] = 90;
// bram[34758] = 72;
// bram[34759] = 55;
// bram[34760] = 40;
// bram[34761] = 26;
// bram[34762] = 16;
// bram[34763] = 7;
// bram[34764] = 2;
// bram[34765] = 0;
// bram[34766] = 0;
// bram[34767] = 4;
// bram[34768] = 10;
// bram[34769] = 19;
// bram[34770] = 31;
// bram[34771] = 45;
// bram[34772] = 61;
// bram[34773] = 79;
// bram[34774] = 97;
// bram[34775] = 117;
// bram[34776] = 136;
// bram[34777] = 155;
// bram[34778] = 174;
// bram[34779] = 191;
// bram[34780] = 207;
// bram[34781] = 221;
// bram[34782] = 233;
// bram[34783] = 243;
// bram[34784] = 249;
// bram[34785] = 253;
// bram[34786] = 253;
// bram[34787] = 251;
// bram[34788] = 246;
// bram[34789] = 238;
// bram[34790] = 227;
// bram[34791] = 214;
// bram[34792] = 199;
// bram[34793] = 182;
// bram[34794] = 163;
// bram[34795] = 144;
// bram[34796] = 125;
// bram[34797] = 105;
// bram[34798] = 86;
// bram[34799] = 68;
// bram[34800] = 52;
// bram[34801] = 37;
// bram[34802] = 24;
// bram[34803] = 14;
// bram[34804] = 6;
// bram[34805] = 1;
// bram[34806] = 0;
// bram[34807] = 1;
// bram[34808] = 5;
// bram[34809] = 12;
// bram[34810] = 21;
// bram[34811] = 34;
// bram[34812] = 48;
// bram[34813] = 64;
// bram[34814] = 82;
// bram[34815] = 101;
// bram[34816] = 120;
// bram[34817] = 140;
// bram[34818] = 159;
// bram[34819] = 177;
// bram[34820] = 195;
// bram[34821] = 210;
// bram[34822] = 224;
// bram[34823] = 235;
// bram[34824] = 244;
// bram[34825] = 250;
// bram[34826] = 253;
// bram[34827] = 253;
// bram[34828] = 250;
// bram[34829] = 244;
// bram[34830] = 236;
// bram[34831] = 225;
// bram[34832] = 211;
// bram[34833] = 196;
// bram[34834] = 178;
// bram[34835] = 160;
// bram[34836] = 141;
// bram[34837] = 121;
// bram[34838] = 102;
// bram[34839] = 83;
// bram[34840] = 65;
// bram[34841] = 49;
// bram[34842] = 34;
// bram[34843] = 22;
// bram[34844] = 12;
// bram[34845] = 5;
// bram[34846] = 1;
// bram[34847] = 0;
// bram[34848] = 1;
// bram[34849] = 6;
// bram[34850] = 13;
// bram[34851] = 24;
// bram[34852] = 36;
// bram[34853] = 51;
// bram[34854] = 67;
// bram[34855] = 85;
// bram[34856] = 104;
// bram[34857] = 124;
// bram[34858] = 143;
// bram[34859] = 162;
// bram[34860] = 181;
// bram[34861] = 198;
// bram[34862] = 213;
// bram[34863] = 226;
// bram[34864] = 237;
// bram[34865] = 245;
// bram[34866] = 251;
// bram[34867] = 253;
// bram[34868] = 253;
// bram[34869] = 249;
// bram[34870] = 243;
// bram[34871] = 234;
// bram[34872] = 222;
// bram[34873] = 208;
// bram[34874] = 193;
// bram[34875] = 175;
// bram[34876] = 157;
// bram[34877] = 137;
// bram[34878] = 118;
// bram[34879] = 98;
// bram[34880] = 80;
// bram[34881] = 62;
// bram[34882] = 46;
// bram[34883] = 32;
// bram[34884] = 20;
// bram[34885] = 11;
// bram[34886] = 4;
// bram[34887] = 0;
// bram[34888] = 0;
// bram[34889] = 2;
// bram[34890] = 7;
// bram[34891] = 15;
// bram[34892] = 26;
// bram[34893] = 39;
// bram[34894] = 54;
// bram[34895] = 71;
// bram[34896] = 89;
// bram[34897] = 108;
// bram[34898] = 127;
// bram[34899] = 147;
// bram[34900] = 166;
// bram[34901] = 184;
// bram[34902] = 201;
// bram[34903] = 215;
// bram[34904] = 228;
// bram[34905] = 239;
// bram[34906] = 247;
// bram[34907] = 251;
// bram[34908] = 253;
// bram[34909] = 252;
// bram[34910] = 248;
// bram[34911] = 242;
// bram[34912] = 232;
// bram[34913] = 220;
// bram[34914] = 206;
// bram[34915] = 189;
// bram[34916] = 172;
// bram[34917] = 153;
// bram[34918] = 134;
// bram[34919] = 114;
// bram[34920] = 95;
// bram[34921] = 76;
// bram[34922] = 59;
// bram[34923] = 43;
// bram[34924] = 30;
// bram[34925] = 18;
// bram[34926] = 9;
// bram[34927] = 3;
// bram[34928] = 0;
// bram[34929] = 0;
// bram[34930] = 3;
// bram[34931] = 8;
// bram[34932] = 17;
// bram[34933] = 28;
// bram[34934] = 41;
// bram[34935] = 57;
// bram[34936] = 74;
// bram[34937] = 92;
// bram[34938] = 111;
// bram[34939] = 131;
// bram[34940] = 150;
// bram[34941] = 169;
// bram[34942] = 187;
// bram[34943] = 203;
// bram[34944] = 218;
// bram[34945] = 230;
// bram[34946] = 240;
// bram[34947] = 248;
// bram[34948] = 252;
// bram[34949] = 253;
// bram[34950] = 252;
// bram[34951] = 247;
// bram[34952] = 240;
// bram[34953] = 230;
// bram[34954] = 217;
// bram[34955] = 203;
// bram[34956] = 186;
// bram[34957] = 168;
// bram[34958] = 150;
// bram[34959] = 130;
// bram[34960] = 111;
// bram[34961] = 91;
// bram[34962] = 73;
// bram[34963] = 56;
// bram[34964] = 41;
// bram[34965] = 27;
// bram[34966] = 16;
// bram[34967] = 8;
// bram[34968] = 2;
// bram[34969] = 0;
// bram[34970] = 0;
// bram[34971] = 3;
// bram[34972] = 10;
// bram[34973] = 19;
// bram[34974] = 30;
// bram[34975] = 44;
// bram[34976] = 60;
// bram[34977] = 77;
// bram[34978] = 96;
// bram[34979] = 115;
// bram[34980] = 134;
// bram[34981] = 154;
// bram[34982] = 173;
// bram[34983] = 190;
// bram[34984] = 206;
// bram[34985] = 220;
// bram[34986] = 232;
// bram[34987] = 242;
// bram[34988] = 249;
// bram[34989] = 253;
// bram[34990] = 253;
// bram[34991] = 251;
// bram[34992] = 246;
// bram[34993] = 238;
// bram[34994] = 228;
// bram[34995] = 215;
// bram[34996] = 200;
// bram[34997] = 183;
// bram[34998] = 165;
// bram[34999] = 146;
// bram[35000] = 127;
// bram[35001] = 107;
// bram[35002] = 88;
// bram[35003] = 70;
// bram[35004] = 53;
// bram[35005] = 38;
// bram[35006] = 25;
// bram[35007] = 15;
// bram[35008] = 7;
// bram[35009] = 2;
// bram[35010] = 0;
// bram[35011] = 0;
// bram[35012] = 4;
// bram[35013] = 11;
// bram[35014] = 21;
// bram[35015] = 33;
// bram[35016] = 47;
// bram[35017] = 63;
// bram[35018] = 80;
// bram[35019] = 99;
// bram[35020] = 119;
// bram[35021] = 138;
// bram[35022] = 157;
// bram[35023] = 176;
// bram[35024] = 193;
// bram[35025] = 209;
// bram[35026] = 223;
// bram[35027] = 234;
// bram[35028] = 243;
// bram[35029] = 250;
// bram[35030] = 253;
// bram[35031] = 253;
// bram[35032] = 251;
// bram[35033] = 245;
// bram[35034] = 237;
// bram[35035] = 226;
// bram[35036] = 212;
// bram[35037] = 197;
// bram[35038] = 180;
// bram[35039] = 162;
// bram[35040] = 142;
// bram[35041] = 123;
// bram[35042] = 103;
// bram[35043] = 85;
// bram[35044] = 67;
// bram[35045] = 50;
// bram[35046] = 36;
// bram[35047] = 23;
// bram[35048] = 13;
// bram[35049] = 6;
// bram[35050] = 1;
// bram[35051] = 0;
// bram[35052] = 1;
// bram[35053] = 5;
// bram[35054] = 13;
// bram[35055] = 23;
// bram[35056] = 35;
// bram[35057] = 50;
// bram[35058] = 66;
// bram[35059] = 84;
// bram[35060] = 103;
// bram[35061] = 122;
// bram[35062] = 142;
// bram[35063] = 161;
// bram[35064] = 179;
// bram[35065] = 196;
// bram[35066] = 212;
// bram[35067] = 225;
// bram[35068] = 236;
// bram[35069] = 245;
// bram[35070] = 250;
// bram[35071] = 253;
// bram[35072] = 253;
// bram[35073] = 250;
// bram[35074] = 244;
// bram[35075] = 235;
// bram[35076] = 223;
// bram[35077] = 210;
// bram[35078] = 194;
// bram[35079] = 177;
// bram[35080] = 158;
// bram[35081] = 139;
// bram[35082] = 119;
// bram[35083] = 100;
// bram[35084] = 81;
// bram[35085] = 64;
// bram[35086] = 47;
// bram[35087] = 33;
// bram[35088] = 21;
// bram[35089] = 11;
// bram[35090] = 5;
// bram[35091] = 1;
// bram[35092] = 0;
// bram[35093] = 2;
// bram[35094] = 6;
// bram[35095] = 14;
// bram[35096] = 25;
// bram[35097] = 38;
// bram[35098] = 52;
// bram[35099] = 69;
// bram[35100] = 87;
// bram[35101] = 106;
// bram[35102] = 126;
// bram[35103] = 145;
// bram[35104] = 164;
// bram[35105] = 182;
// bram[35106] = 199;
// bram[35107] = 214;
// bram[35108] = 227;
// bram[35109] = 238;
// bram[35110] = 246;
// bram[35111] = 251;
// bram[35112] = 253;
// bram[35113] = 253;
// bram[35114] = 249;
// bram[35115] = 242;
// bram[35116] = 233;
// bram[35117] = 221;
// bram[35118] = 207;
// bram[35119] = 191;
// bram[35120] = 173;
// bram[35121] = 155;
// bram[35122] = 135;
// bram[35123] = 116;
// bram[35124] = 96;
// bram[35125] = 78;
// bram[35126] = 60;
// bram[35127] = 45;
// bram[35128] = 31;
// bram[35129] = 19;
// bram[35130] = 10;
// bram[35131] = 4;
// bram[35132] = 0;
// bram[35133] = 0;
// bram[35134] = 2;
// bram[35135] = 8;
// bram[35136] = 16;
// bram[35137] = 27;
// bram[35138] = 40;
// bram[35139] = 55;
// bram[35140] = 72;
// bram[35141] = 91;
// bram[35142] = 110;
// bram[35143] = 129;
// bram[35144] = 149;
// bram[35145] = 168;
// bram[35146] = 186;
// bram[35147] = 202;
// bram[35148] = 217;
// bram[35149] = 229;
// bram[35150] = 240;
// bram[35151] = 247;
// bram[35152] = 252;
// bram[35153] = 253;
// bram[35154] = 252;
// bram[35155] = 248;
// bram[35156] = 241;
// bram[35157] = 231;
// bram[35158] = 219;
// bram[35159] = 204;
// bram[35160] = 188;
// bram[35161] = 170;
// bram[35162] = 151;
// bram[35163] = 132;
// bram[35164] = 112;
// bram[35165] = 93;
// bram[35166] = 75;
// bram[35167] = 57;
// bram[35168] = 42;
// bram[35169] = 28;
// bram[35170] = 17;
// bram[35171] = 9;
// bram[35172] = 3;
// bram[35173] = 0;
// bram[35174] = 0;
// bram[35175] = 3;
// bram[35176] = 9;
// bram[35177] = 18;
// bram[35178] = 29;
// bram[35179] = 43;
// bram[35180] = 58;
// bram[35181] = 76;
// bram[35182] = 94;
// bram[35183] = 113;
// bram[35184] = 133;
// bram[35185] = 152;
// bram[35186] = 171;
// bram[35187] = 189;
// bram[35188] = 205;
// bram[35189] = 219;
// bram[35190] = 232;
// bram[35191] = 241;
// bram[35192] = 248;
// bram[35193] = 252;
// bram[35194] = 253;
// bram[35195] = 252;
// bram[35196] = 247;
// bram[35197] = 239;
// bram[35198] = 229;
// bram[35199] = 216;
// bram[35200] = 201;
// bram[35201] = 185;
// bram[35202] = 167;
// bram[35203] = 148;
// bram[35204] = 128;
// bram[35205] = 109;
// bram[35206] = 90;
// bram[35207] = 71;
// bram[35208] = 54;
// bram[35209] = 39;
// bram[35210] = 26;
// bram[35211] = 15;
// bram[35212] = 7;
// bram[35213] = 2;
// bram[35214] = 0;
// bram[35215] = 0;
// bram[35216] = 4;
// bram[35217] = 10;
// bram[35218] = 20;
// bram[35219] = 32;
// bram[35220] = 46;
// bram[35221] = 62;
// bram[35222] = 79;
// bram[35223] = 98;
// bram[35224] = 117;
// bram[35225] = 136;
// bram[35226] = 156;
// bram[35227] = 174;
// bram[35228] = 192;
// bram[35229] = 208;
// bram[35230] = 222;
// bram[35231] = 234;
// bram[35232] = 243;
// bram[35233] = 249;
// bram[35234] = 253;
// bram[35235] = 253;
// bram[35236] = 251;
// bram[35237] = 246;
// bram[35238] = 237;
// bram[35239] = 227;
// bram[35240] = 213;
// bram[35241] = 198;
// bram[35242] = 181;
// bram[35243] = 163;
// bram[35244] = 144;
// bram[35245] = 125;
// bram[35246] = 105;
// bram[35247] = 86;
// bram[35248] = 68;
// bram[35249] = 52;
// bram[35250] = 37;
// bram[35251] = 24;
// bram[35252] = 14;
// bram[35253] = 6;
// bram[35254] = 1;
// bram[35255] = 0;
// bram[35256] = 1;
// bram[35257] = 5;
// bram[35258] = 12;
// bram[35259] = 22;
// bram[35260] = 34;
// bram[35261] = 48;
// bram[35262] = 65;
// bram[35263] = 82;
// bram[35264] = 101;
// bram[35265] = 121;
// bram[35266] = 140;
// bram[35267] = 159;
// bram[35268] = 178;
// bram[35269] = 195;
// bram[35270] = 210;
// bram[35271] = 224;
// bram[35272] = 235;
// bram[35273] = 244;
// bram[35274] = 250;
// bram[35275] = 253;
// bram[35276] = 253;
// bram[35277] = 250;
// bram[35278] = 244;
// bram[35279] = 236;
// bram[35280] = 224;
// bram[35281] = 211;
// bram[35282] = 195;
// bram[35283] = 178;
// bram[35284] = 160;
// bram[35285] = 140;
// bram[35286] = 121;
// bram[35287] = 102;
// bram[35288] = 83;
// bram[35289] = 65;
// bram[35290] = 49;
// bram[35291] = 34;
// bram[35292] = 22;
// bram[35293] = 12;
// bram[35294] = 5;
// bram[35295] = 1;
// bram[35296] = 0;
// bram[35297] = 1;
// bram[35298] = 6;
// bram[35299] = 14;
// bram[35300] = 24;
// bram[35301] = 36;
// bram[35302] = 51;
// bram[35303] = 68;
// bram[35304] = 86;
// bram[35305] = 105;
// bram[35306] = 124;
// bram[35307] = 144;
// bram[35308] = 163;
// bram[35309] = 181;
// bram[35310] = 198;
// bram[35311] = 213;
// bram[35312] = 226;
// bram[35313] = 237;
// bram[35314] = 245;
// bram[35315] = 251;
// bram[35316] = 253;
// bram[35317] = 253;
// bram[35318] = 249;
// bram[35319] = 243;
// bram[35320] = 234;
// bram[35321] = 222;
// bram[35322] = 208;
// bram[35323] = 192;
// bram[35324] = 175;
// bram[35325] = 156;
// bram[35326] = 137;
// bram[35327] = 117;
// bram[35328] = 98;
// bram[35329] = 79;
// bram[35330] = 62;
// bram[35331] = 46;
// bram[35332] = 32;
// bram[35333] = 20;
// bram[35334] = 11;
// bram[35335] = 4;
// bram[35336] = 0;
// bram[35337] = 0;
// bram[35338] = 2;
// bram[35339] = 7;
// bram[35340] = 15;
// bram[35341] = 26;
// bram[35342] = 39;
// bram[35343] = 54;
// bram[35344] = 71;
// bram[35345] = 89;
// bram[35346] = 108;
// bram[35347] = 128;
// bram[35348] = 147;
// bram[35349] = 166;
// bram[35350] = 184;
// bram[35351] = 201;
// bram[35352] = 216;
// bram[35353] = 229;
// bram[35354] = 239;
// bram[35355] = 247;
// bram[35356] = 252;
// bram[35357] = 253;
// bram[35358] = 252;
// bram[35359] = 248;
// bram[35360] = 241;
// bram[35361] = 232;
// bram[35362] = 220;
// bram[35363] = 205;
// bram[35364] = 189;
// bram[35365] = 171;
// bram[35366] = 153;
// bram[35367] = 133;
// bram[35368] = 114;
// bram[35369] = 95;
// bram[35370] = 76;
// bram[35371] = 59;
// bram[35372] = 43;
// bram[35373] = 29;
// bram[35374] = 18;
// bram[35375] = 9;
// bram[35376] = 3;
// bram[35377] = 0;
// bram[35378] = 0;
// bram[35379] = 3;
// bram[35380] = 8;
// bram[35381] = 17;
// bram[35382] = 28;
// bram[35383] = 42;
// bram[35384] = 57;
// bram[35385] = 74;
// bram[35386] = 93;
// bram[35387] = 112;
// bram[35388] = 131;
// bram[35389] = 151;
// bram[35390] = 170;
// bram[35391] = 187;
// bram[35392] = 204;
// bram[35393] = 218;
// bram[35394] = 231;
// bram[35395] = 241;
// bram[35396] = 248;
// bram[35397] = 252;
// bram[35398] = 253;
// bram[35399] = 252;
// bram[35400] = 247;
// bram[35401] = 240;
// bram[35402] = 230;
// bram[35403] = 217;
// bram[35404] = 202;
// bram[35405] = 186;
// bram[35406] = 168;
// bram[35407] = 149;
// bram[35408] = 130;
// bram[35409] = 110;
// bram[35410] = 91;
// bram[35411] = 73;
// bram[35412] = 56;
// bram[35413] = 40;
// bram[35414] = 27;
// bram[35415] = 16;
// bram[35416] = 8;
// bram[35417] = 2;
// bram[35418] = 0;
// bram[35419] = 0;
// bram[35420] = 3;
// bram[35421] = 10;
// bram[35422] = 19;
// bram[35423] = 30;
// bram[35424] = 44;
// bram[35425] = 60;
// bram[35426] = 78;
// bram[35427] = 96;
// bram[35428] = 115;
// bram[35429] = 135;
// bram[35430] = 154;
// bram[35431] = 173;
// bram[35432] = 190;
// bram[35433] = 207;
// bram[35434] = 221;
// bram[35435] = 233;
// bram[35436] = 242;
// bram[35437] = 249;
// bram[35438] = 253;
// bram[35439] = 253;
// bram[35440] = 251;
// bram[35441] = 246;
// bram[35442] = 238;
// bram[35443] = 228;
// bram[35444] = 215;
// bram[35445] = 200;
// bram[35446] = 183;
// bram[35447] = 165;
// bram[35448] = 146;
// bram[35449] = 126;
// bram[35450] = 107;
// bram[35451] = 88;
// bram[35452] = 70;
// bram[35453] = 53;
// bram[35454] = 38;
// bram[35455] = 25;
// bram[35456] = 14;
// bram[35457] = 7;
// bram[35458] = 2;
// bram[35459] = 0;
// bram[35460] = 1;
// bram[35461] = 4;
// bram[35462] = 11;
// bram[35463] = 21;
// bram[35464] = 33;
// bram[35465] = 47;
// bram[35466] = 63;
// bram[35467] = 81;
// bram[35468] = 100;
// bram[35469] = 119;
// bram[35470] = 138;
// bram[35471] = 158;
// bram[35472] = 176;
// bram[35473] = 194;
// bram[35474] = 209;
// bram[35475] = 223;
// bram[35476] = 235;
// bram[35477] = 244;
// bram[35478] = 250;
// bram[35479] = 253;
// bram[35480] = 253;
// bram[35481] = 251;
// bram[35482] = 245;
// bram[35483] = 236;
// bram[35484] = 225;
// bram[35485] = 212;
// bram[35486] = 197;
// bram[35487] = 179;
// bram[35488] = 161;
// bram[35489] = 142;
// bram[35490] = 123;
// bram[35491] = 103;
// bram[35492] = 84;
// bram[35493] = 66;
// bram[35494] = 50;
// bram[35495] = 35;
// bram[35496] = 23;
// bram[35497] = 13;
// bram[35498] = 5;
// bram[35499] = 1;
// bram[35500] = 0;
// bram[35501] = 1;
// bram[35502] = 5;
// bram[35503] = 13;
// bram[35504] = 23;
// bram[35505] = 35;
// bram[35506] = 50;
// bram[35507] = 66;
// bram[35508] = 84;
// bram[35509] = 103;
// bram[35510] = 123;
// bram[35511] = 142;
// bram[35512] = 161;
// bram[35513] = 179;
// bram[35514] = 197;
// bram[35515] = 212;
// bram[35516] = 225;
// bram[35517] = 236;
// bram[35518] = 245;
// bram[35519] = 251;
// bram[35520] = 253;
// bram[35521] = 253;
// bram[35522] = 250;
// bram[35523] = 244;
// bram[35524] = 235;
// bram[35525] = 223;
// bram[35526] = 209;
// bram[35527] = 194;
// bram[35528] = 176;
// bram[35529] = 158;
// bram[35530] = 138;
// bram[35531] = 119;
// bram[35532] = 100;
// bram[35533] = 81;
// bram[35534] = 63;
// bram[35535] = 47;
// bram[35536] = 33;
// bram[35537] = 21;
// bram[35538] = 11;
// bram[35539] = 4;
// bram[35540] = 1;
// bram[35541] = 0;
// bram[35542] = 2;
// bram[35543] = 7;
// bram[35544] = 14;
// bram[35545] = 25;
// bram[35546] = 38;
// bram[35547] = 53;
// bram[35548] = 70;
// bram[35549] = 88;
// bram[35550] = 107;
// bram[35551] = 126;
// bram[35552] = 146;
// bram[35553] = 165;
// bram[35554] = 183;
// bram[35555] = 200;
// bram[35556] = 215;
// bram[35557] = 228;
// bram[35558] = 238;
// bram[35559] = 246;
// bram[35560] = 251;
// bram[35561] = 253;
// bram[35562] = 253;
// bram[35563] = 249;
// bram[35564] = 242;
// bram[35565] = 233;
// bram[35566] = 221;
// bram[35567] = 207;
// bram[35568] = 190;
// bram[35569] = 173;
// bram[35570] = 154;
// bram[35571] = 135;
// bram[35572] = 115;
// bram[35573] = 96;
// bram[35574] = 78;
// bram[35575] = 60;
// bram[35576] = 44;
// bram[35577] = 30;
// bram[35578] = 19;
// bram[35579] = 10;
// bram[35580] = 3;
// bram[35581] = 0;
// bram[35582] = 0;
// bram[35583] = 2;
// bram[35584] = 8;
// bram[35585] = 16;
// bram[35586] = 27;
// bram[35587] = 40;
// bram[35588] = 56;
// bram[35589] = 73;
// bram[35590] = 91;
// bram[35591] = 110;
// bram[35592] = 130;
// bram[35593] = 149;
// bram[35594] = 168;
// bram[35595] = 186;
// bram[35596] = 202;
// bram[35597] = 217;
// bram[35598] = 230;
// bram[35599] = 240;
// bram[35600] = 247;
// bram[35601] = 252;
// bram[35602] = 253;
// bram[35603] = 252;
// bram[35604] = 248;
// bram[35605] = 241;
// bram[35606] = 231;
// bram[35607] = 218;
// bram[35608] = 204;
// bram[35609] = 187;
// bram[35610] = 170;
// bram[35611] = 151;
// bram[35612] = 131;
// bram[35613] = 112;
// bram[35614] = 93;
// bram[35615] = 74;
// bram[35616] = 57;
// bram[35617] = 42;
// bram[35618] = 28;
// bram[35619] = 17;
// bram[35620] = 8;
// bram[35621] = 3;
// bram[35622] = 0;
// bram[35623] = 0;
// bram[35624] = 3;
// bram[35625] = 9;
// bram[35626] = 18;
// bram[35627] = 29;
// bram[35628] = 43;
// bram[35629] = 59;
// bram[35630] = 76;
// bram[35631] = 95;
// bram[35632] = 114;
// bram[35633] = 133;
// bram[35634] = 153;
// bram[35635] = 171;
// bram[35636] = 189;
// bram[35637] = 205;
// bram[35638] = 220;
// bram[35639] = 232;
// bram[35640] = 241;
// bram[35641] = 248;
// bram[35642] = 252;
// bram[35643] = 253;
// bram[35644] = 252;
// bram[35645] = 247;
// bram[35646] = 239;
// bram[35647] = 229;
// bram[35648] = 216;
// bram[35649] = 201;
// bram[35650] = 184;
// bram[35651] = 166;
// bram[35652] = 147;
// bram[35653] = 128;
// bram[35654] = 108;
// bram[35655] = 89;
// bram[35656] = 71;
// bram[35657] = 54;
// bram[35658] = 39;
// bram[35659] = 26;
// bram[35660] = 15;
// bram[35661] = 7;
// bram[35662] = 2;
// bram[35663] = 0;
// bram[35664] = 0;
// bram[35665] = 4;
// bram[35666] = 11;
// bram[35667] = 20;
// bram[35668] = 32;
// bram[35669] = 46;
// bram[35670] = 62;
// bram[35671] = 79;
// bram[35672] = 98;
// bram[35673] = 117;
// bram[35674] = 137;
// bram[35675] = 156;
// bram[35676] = 175;
// bram[35677] = 192;
// bram[35678] = 208;
// bram[35679] = 222;
// bram[35680] = 234;
// bram[35681] = 243;
// bram[35682] = 249;
// bram[35683] = 253;
// bram[35684] = 253;
// bram[35685] = 251;
// bram[35686] = 245;
// bram[35687] = 237;
// bram[35688] = 226;
// bram[35689] = 213;
// bram[35690] = 198;
// bram[35691] = 181;
// bram[35692] = 163;
// bram[35693] = 144;
// bram[35694] = 124;
// bram[35695] = 105;
// bram[35696] = 86;
// bram[35697] = 68;
// bram[35698] = 51;
// bram[35699] = 36;
// bram[35700] = 24;
// bram[35701] = 14;
// bram[35702] = 6;
// bram[35703] = 1;
// bram[35704] = 0;
// bram[35705] = 1;
// bram[35706] = 5;
// bram[35707] = 12;
// bram[35708] = 22;
// bram[35709] = 34;
// bram[35710] = 49;
// bram[35711] = 65;
// bram[35712] = 83;
// bram[35713] = 102;
// bram[35714] = 121;
// bram[35715] = 140;
// bram[35716] = 160;
// bram[35717] = 178;
// bram[35718] = 195;
// bram[35719] = 211;
// bram[35720] = 224;
// bram[35721] = 236;
// bram[35722] = 244;
// bram[35723] = 250;
// bram[35724] = 253;
// bram[35725] = 253;
// bram[35726] = 250;
// bram[35727] = 244;
// bram[35728] = 235;
// bram[35729] = 224;
// bram[35730] = 210;
// bram[35731] = 195;
// bram[35732] = 178;
// bram[35733] = 159;
// bram[35734] = 140;
// bram[35735] = 121;
// bram[35736] = 101;
// bram[35737] = 82;
// bram[35738] = 65;
// bram[35739] = 48;
// bram[35740] = 34;
// bram[35741] = 22;
// bram[35742] = 12;
// bram[35743] = 5;
// bram[35744] = 1;
// bram[35745] = 0;
// bram[35746] = 1;
// bram[35747] = 6;
// bram[35748] = 14;
// bram[35749] = 24;
// bram[35750] = 37;
// bram[35751] = 52;
// bram[35752] = 68;
// bram[35753] = 86;
// bram[35754] = 105;
// bram[35755] = 125;
// bram[35756] = 144;
// bram[35757] = 163;
// bram[35758] = 181;
// bram[35759] = 198;
// bram[35760] = 213;
// bram[35761] = 227;
// bram[35762] = 237;
// bram[35763] = 246;
// bram[35764] = 251;
// bram[35765] = 253;
// bram[35766] = 253;
// bram[35767] = 249;
// bram[35768] = 243;
// bram[35769] = 234;
// bram[35770] = 222;
// bram[35771] = 208;
// bram[35772] = 192;
// bram[35773] = 174;
// bram[35774] = 156;
// bram[35775] = 136;
// bram[35776] = 117;
// bram[35777] = 98;
// bram[35778] = 79;
// bram[35779] = 62;
// bram[35780] = 46;
// bram[35781] = 32;
// bram[35782] = 20;
// bram[35783] = 10;
// bram[35784] = 4;
// bram[35785] = 0;
// bram[35786] = 0;
// bram[35787] = 2;
// bram[35788] = 7;
// bram[35789] = 15;
// bram[35790] = 26;
// bram[35791] = 39;
// bram[35792] = 54;
// bram[35793] = 71;
// bram[35794] = 90;
// bram[35795] = 109;
// bram[35796] = 128;
// bram[35797] = 148;
// bram[35798] = 167;
// bram[35799] = 185;
// bram[35800] = 201;
// bram[35801] = 216;
// bram[35802] = 229;
// bram[35803] = 239;
// bram[35804] = 247;
// bram[35805] = 252;
// bram[35806] = 253;
// bram[35807] = 252;
// bram[35808] = 248;
// bram[35809] = 241;
// bram[35810] = 232;
// bram[35811] = 219;
// bram[35812] = 205;
// bram[35813] = 189;
// bram[35814] = 171;
// bram[35815] = 152;
// bram[35816] = 133;
// bram[35817] = 113;
// bram[35818] = 94;
// bram[35819] = 76;
// bram[35820] = 58;
// bram[35821] = 43;
// bram[35822] = 29;
// bram[35823] = 18;
// bram[35824] = 9;
// bram[35825] = 3;
// bram[35826] = 0;
// bram[35827] = 0;
// bram[35828] = 3;
// bram[35829] = 9;
// bram[35830] = 17;
// bram[35831] = 28;
// bram[35832] = 42;
// bram[35833] = 57;
// bram[35834] = 75;
// bram[35835] = 93;
// bram[35836] = 112;
// bram[35837] = 132;
// bram[35838] = 151;
// bram[35839] = 170;
// bram[35840] = 188;
// bram[35841] = 204;
// bram[35842] = 219;
// bram[35843] = 231;
// bram[35844] = 241;
// bram[35845] = 248;
// bram[35846] = 252;
// bram[35847] = 253;
// bram[35848] = 252;
// bram[35849] = 247;
// bram[35850] = 240;
// bram[35851] = 229;
// bram[35852] = 217;
// bram[35853] = 202;
// bram[35854] = 186;
// bram[35855] = 168;
// bram[35856] = 149;
// bram[35857] = 129;
// bram[35858] = 110;
// bram[35859] = 91;
// bram[35860] = 72;
// bram[35861] = 55;
// bram[35862] = 40;
// bram[35863] = 27;
// bram[35864] = 16;
// bram[35865] = 8;
// bram[35866] = 2;
// bram[35867] = 0;
// bram[35868] = 0;
// bram[35869] = 4;
// bram[35870] = 10;
// bram[35871] = 19;
// bram[35872] = 31;
// bram[35873] = 45;
// bram[35874] = 60;
// bram[35875] = 78;
// bram[35876] = 96;
// bram[35877] = 116;
// bram[35878] = 135;
// bram[35879] = 155;
// bram[35880] = 173;
// bram[35881] = 191;
// bram[35882] = 207;
// bram[35883] = 221;
// bram[35884] = 233;
// bram[35885] = 242;
// bram[35886] = 249;
// bram[35887] = 253;
// bram[35888] = 253;
// bram[35889] = 251;
// bram[35890] = 246;
// bram[35891] = 238;
// bram[35892] = 227;
// bram[35893] = 214;
// bram[35894] = 199;
// bram[35895] = 182;
// bram[35896] = 164;
// bram[35897] = 145;
// bram[35898] = 126;
// bram[35899] = 106;
// bram[35900] = 87;
// bram[35901] = 69;
// bram[35902] = 52;
// bram[35903] = 38;
// bram[35904] = 25;
// bram[35905] = 14;
// bram[35906] = 6;
// bram[35907] = 2;
// bram[35908] = 0;
// bram[35909] = 1;
// bram[35910] = 5;
// bram[35911] = 11;
// bram[35912] = 21;
// bram[35913] = 33;
// bram[35914] = 47;
// bram[35915] = 64;
// bram[35916] = 81;
// bram[35917] = 100;
// bram[35918] = 119;
// bram[35919] = 139;
// bram[35920] = 158;
// bram[35921] = 177;
// bram[35922] = 194;
// bram[35923] = 210;
// bram[35924] = 223;
// bram[35925] = 235;
// bram[35926] = 244;
// bram[35927] = 250;
// bram[35928] = 253;
// bram[35929] = 253;
// bram[35930] = 250;
// bram[35931] = 245;
// bram[35932] = 236;
// bram[35933] = 225;
// bram[35934] = 212;
// bram[35935] = 196;
// bram[35936] = 179;
// bram[35937] = 161;
// bram[35938] = 142;
// bram[35939] = 122;
// bram[35940] = 103;
// bram[35941] = 84;
// bram[35942] = 66;
// bram[35943] = 50;
// bram[35944] = 35;
// bram[35945] = 23;
// bram[35946] = 13;
// bram[35947] = 5;
// bram[35948] = 1;
// bram[35949] = 0;
// bram[35950] = 1;
// bram[35951] = 6;
// bram[35952] = 13;
// bram[35953] = 23;
// bram[35954] = 36;
// bram[35955] = 50;
// bram[35956] = 67;
// bram[35957] = 85;
// bram[35958] = 103;
// bram[35959] = 123;
// bram[35960] = 142;
// bram[35961] = 162;
// bram[35962] = 180;
// bram[35963] = 197;
// bram[35964] = 212;
// bram[35965] = 226;
// bram[35966] = 237;
// bram[35967] = 245;
// bram[35968] = 251;
// bram[35969] = 253;
// bram[35970] = 253;
// bram[35971] = 250;
// bram[35972] = 243;
// bram[35973] = 234;
// bram[35974] = 223;
// bram[35975] = 209;
// bram[35976] = 193;
// bram[35977] = 176;
// bram[35978] = 157;
// bram[35979] = 138;
// bram[35980] = 119;
// bram[35981] = 99;
// bram[35982] = 80;
// bram[35983] = 63;
// bram[35984] = 47;
// bram[35985] = 33;
// bram[35986] = 21;
// bram[35987] = 11;
// bram[35988] = 4;
// bram[35989] = 0;
// bram[35990] = 0;
// bram[35991] = 2;
// bram[35992] = 7;
// bram[35993] = 15;
// bram[35994] = 25;
// bram[35995] = 38;
// bram[35996] = 53;
// bram[35997] = 70;
// bram[35998] = 88;
// bram[35999] = 107;
// bram[36000] = 126;
// bram[36001] = 146;
// bram[36002] = 165;
// bram[36003] = 183;
// bram[36004] = 200;
// bram[36005] = 215;
// bram[36006] = 228;
// bram[36007] = 238;
// bram[36008] = 246;
// bram[36009] = 251;
// bram[36010] = 253;
// bram[36011] = 253;
// bram[36012] = 249;
// bram[36013] = 242;
// bram[36014] = 232;
// bram[36015] = 220;
// bram[36016] = 206;
// bram[36017] = 190;
// bram[36018] = 173;
// bram[36019] = 154;
// bram[36020] = 134;
// bram[36021] = 115;
// bram[36022] = 96;
// bram[36023] = 77;
// bram[36024] = 60;
// bram[36025] = 44;
// bram[36026] = 30;
// bram[36027] = 19;
// bram[36028] = 10;
// bram[36029] = 3;
// bram[36030] = 0;
// bram[36031] = 0;
// bram[36032] = 2;
// bram[36033] = 8;
// bram[36034] = 16;
// bram[36035] = 27;
// bram[36036] = 41;
// bram[36037] = 56;
// bram[36038] = 73;
// bram[36039] = 91;
// bram[36040] = 111;
// bram[36041] = 130;
// bram[36042] = 150;
// bram[36043] = 168;
// bram[36044] = 186;
// bram[36045] = 203;
// bram[36046] = 217;
// bram[36047] = 230;
// bram[36048] = 240;
// bram[36049] = 247;
// bram[36050] = 252;
// bram[36051] = 253;
// bram[36052] = 252;
// bram[36053] = 248;
// bram[36054] = 240;
// bram[36055] = 230;
// bram[36056] = 218;
// bram[36057] = 203;
// bram[36058] = 187;
// bram[36059] = 169;
// bram[36060] = 150;
// bram[36061] = 131;
// bram[36062] = 111;
// bram[36063] = 92;
// bram[36064] = 74;
// bram[36065] = 57;
// bram[36066] = 41;
// bram[36067] = 28;
// bram[36068] = 17;
// bram[36069] = 8;
// bram[36070] = 3;
// bram[36071] = 0;
// bram[36072] = 0;
// bram[36073] = 3;
// bram[36074] = 9;
// bram[36075] = 18;
// bram[36076] = 30;
// bram[36077] = 43;
// bram[36078] = 59;
// bram[36079] = 76;
// bram[36080] = 95;
// bram[36081] = 114;
// bram[36082] = 134;
// bram[36083] = 153;
// bram[36084] = 172;
// bram[36085] = 189;
// bram[36086] = 206;
// bram[36087] = 220;
// bram[36088] = 232;
// bram[36089] = 242;
// bram[36090] = 248;
// bram[36091] = 252;
// bram[36092] = 253;
// bram[36093] = 251;
// bram[36094] = 247;
// bram[36095] = 239;
// bram[36096] = 228;
// bram[36097] = 215;
// bram[36098] = 201;
// bram[36099] = 184;
// bram[36100] = 166;
// bram[36101] = 147;
// bram[36102] = 127;
// bram[36103] = 108;
// bram[36104] = 89;
// bram[36105] = 71;
// bram[36106] = 54;
// bram[36107] = 39;
// bram[36108] = 26;
// bram[36109] = 15;
// bram[36110] = 7;
// bram[36111] = 2;
// bram[36112] = 0;
// bram[36113] = 0;
// bram[36114] = 4;
// bram[36115] = 11;
// bram[36116] = 20;
// bram[36117] = 32;
// bram[36118] = 46;
// bram[36119] = 62;
// bram[36120] = 80;
// bram[36121] = 98;
// bram[36122] = 118;
// bram[36123] = 137;
// bram[36124] = 157;
// bram[36125] = 175;
// bram[36126] = 193;
// bram[36127] = 208;
// bram[36128] = 222;
// bram[36129] = 234;
// bram[36130] = 243;
// bram[36131] = 249;
// bram[36132] = 253;
// bram[36133] = 253;
// bram[36134] = 251;
// bram[36135] = 245;
// bram[36136] = 237;
// bram[36137] = 226;
// bram[36138] = 213;
// bram[36139] = 198;
// bram[36140] = 181;
// bram[36141] = 162;
// bram[36142] = 143;
// bram[36143] = 124;
// bram[36144] = 104;
// bram[36145] = 85;
// bram[36146] = 67;
// bram[36147] = 51;
// bram[36148] = 36;
// bram[36149] = 24;
// bram[36150] = 13;
// bram[36151] = 6;
// bram[36152] = 1;
// bram[36153] = 0;
// bram[36154] = 1;
// bram[36155] = 5;
// bram[36156] = 12;
// bram[36157] = 22;
// bram[36158] = 34;
// bram[36159] = 49;
// bram[36160] = 65;
// bram[36161] = 83;
// bram[36162] = 102;
// bram[36163] = 121;
// bram[36164] = 141;
// bram[36165] = 160;
// bram[36166] = 178;
// bram[36167] = 196;
// bram[36168] = 211;
// bram[36169] = 225;
// bram[36170] = 236;
// bram[36171] = 244;
// bram[36172] = 250;
// bram[36173] = 253;
// bram[36174] = 253;
// bram[36175] = 250;
// bram[36176] = 244;
// bram[36177] = 235;
// bram[36178] = 224;
// bram[36179] = 210;
// bram[36180] = 195;
// bram[36181] = 177;
// bram[36182] = 159;
// bram[36183] = 140;
// bram[36184] = 120;
// bram[36185] = 101;
// bram[36186] = 82;
// bram[36187] = 64;
// bram[36188] = 48;
// bram[36189] = 34;
// bram[36190] = 21;
// bram[36191] = 12;
// bram[36192] = 5;
// bram[36193] = 1;
// bram[36194] = 0;
// bram[36195] = 1;
// bram[36196] = 6;
// bram[36197] = 14;
// bram[36198] = 24;
// bram[36199] = 37;
// bram[36200] = 52;
// bram[36201] = 68;
// bram[36202] = 86;
// bram[36203] = 105;
// bram[36204] = 125;
// bram[36205] = 144;
// bram[36206] = 163;
// bram[36207] = 182;
// bram[36208] = 199;
// bram[36209] = 214;
// bram[36210] = 227;
// bram[36211] = 238;
// bram[36212] = 246;
// bram[36213] = 251;
// bram[36214] = 253;
// bram[36215] = 253;
// bram[36216] = 249;
// bram[36217] = 243;
// bram[36218] = 233;
// bram[36219] = 221;
// bram[36220] = 207;
// bram[36221] = 191;
// bram[36222] = 174;
// bram[36223] = 155;
// bram[36224] = 136;
// bram[36225] = 117;
// bram[36226] = 97;
// bram[36227] = 79;
// bram[36228] = 61;
// bram[36229] = 45;
// bram[36230] = 31;
// bram[36231] = 19;
// bram[36232] = 10;
// bram[36233] = 4;
// bram[36234] = 0;
// bram[36235] = 0;
// bram[36236] = 2;
// bram[36237] = 7;
// bram[36238] = 16;
// bram[36239] = 26;
// bram[36240] = 40;
// bram[36241] = 55;
// bram[36242] = 72;
// bram[36243] = 90;
// bram[36244] = 109;
// bram[36245] = 128;
// bram[36246] = 148;
// bram[36247] = 167;
// bram[36248] = 185;
// bram[36249] = 201;
// bram[36250] = 216;
// bram[36251] = 229;
// bram[36252] = 239;
// bram[36253] = 247;
// bram[36254] = 252;
// bram[36255] = 253;
// bram[36256] = 252;
// bram[36257] = 248;
// bram[36258] = 241;
// bram[36259] = 231;
// bram[36260] = 219;
// bram[36261] = 205;
// bram[36262] = 188;
// bram[36263] = 171;
// bram[36264] = 152;
// bram[36265] = 132;
// bram[36266] = 113;
// bram[36267] = 94;
// bram[36268] = 75;
// bram[36269] = 58;
// bram[36270] = 43;
// bram[36271] = 29;
// bram[36272] = 18;
// bram[36273] = 9;
// bram[36274] = 3;
// bram[36275] = 0;
// bram[36276] = 0;
// bram[36277] = 3;
// bram[36278] = 9;
// bram[36279] = 17;
// bram[36280] = 29;
// bram[36281] = 42;
// bram[36282] = 58;
// bram[36283] = 75;
// bram[36284] = 93;
// bram[36285] = 113;
// bram[36286] = 132;
// bram[36287] = 151;
// bram[36288] = 170;
// bram[36289] = 188;
// bram[36290] = 204;
// bram[36291] = 219;
// bram[36292] = 231;
// bram[36293] = 241;
// bram[36294] = 248;
// bram[36295] = 252;
// bram[36296] = 253;
// bram[36297] = 252;
// bram[36298] = 247;
// bram[36299] = 239;
// bram[36300] = 229;
// bram[36301] = 217;
// bram[36302] = 202;
// bram[36303] = 185;
// bram[36304] = 167;
// bram[36305] = 148;
// bram[36306] = 129;
// bram[36307] = 109;
// bram[36308] = 90;
// bram[36309] = 72;
// bram[36310] = 55;
// bram[36311] = 40;
// bram[36312] = 27;
// bram[36313] = 16;
// bram[36314] = 8;
// bram[36315] = 2;
// bram[36316] = 0;
// bram[36317] = 0;
// bram[36318] = 4;
// bram[36319] = 10;
// bram[36320] = 19;
// bram[36321] = 31;
// bram[36322] = 45;
// bram[36323] = 61;
// bram[36324] = 78;
// bram[36325] = 97;
// bram[36326] = 116;
// bram[36327] = 136;
// bram[36328] = 155;
// bram[36329] = 174;
// bram[36330] = 191;
// bram[36331] = 207;
// bram[36332] = 221;
// bram[36333] = 233;
// bram[36334] = 242;
// bram[36335] = 249;
// bram[36336] = 253;
// bram[36337] = 253;
// bram[36338] = 251;
// bram[36339] = 246;
// bram[36340] = 238;
// bram[36341] = 227;
// bram[36342] = 214;
// bram[36343] = 199;
// bram[36344] = 182;
// bram[36345] = 164;
// bram[36346] = 145;
// bram[36347] = 125;
// bram[36348] = 106;
// bram[36349] = 87;
// bram[36350] = 69;
// bram[36351] = 52;
// bram[36352] = 37;
// bram[36353] = 24;
// bram[36354] = 14;
// bram[36355] = 6;
// bram[36356] = 1;
// bram[36357] = 0;
// bram[36358] = 1;
// bram[36359] = 5;
// bram[36360] = 12;
// bram[36361] = 21;
// bram[36362] = 33;
// bram[36363] = 48;
// bram[36364] = 64;
// bram[36365] = 82;
// bram[36366] = 100;
// bram[36367] = 120;
// bram[36368] = 139;
// bram[36369] = 158;
// bram[36370] = 177;
// bram[36371] = 194;
// bram[36372] = 210;
// bram[36373] = 224;
// bram[36374] = 235;
// bram[36375] = 244;
// bram[36376] = 250;
// bram[36377] = 253;
// bram[36378] = 253;
// bram[36379] = 250;
// bram[36380] = 245;
// bram[36381] = 236;
// bram[36382] = 225;
// bram[36383] = 211;
// bram[36384] = 196;
// bram[36385] = 179;
// bram[36386] = 160;
// bram[36387] = 141;
// bram[36388] = 122;
// bram[36389] = 102;
// bram[36390] = 83;
// bram[36391] = 66;
// bram[36392] = 49;
// bram[36393] = 35;
// bram[36394] = 22;
// bram[36395] = 12;
// bram[36396] = 5;
// bram[36397] = 1;
// bram[36398] = 0;
// bram[36399] = 1;
// bram[36400] = 6;
// bram[36401] = 13;
// bram[36402] = 23;
// bram[36403] = 36;
// bram[36404] = 51;
// bram[36405] = 67;
// bram[36406] = 85;
// bram[36407] = 104;
// bram[36408] = 123;
// bram[36409] = 143;
// bram[36410] = 162;
// bram[36411] = 180;
// bram[36412] = 197;
// bram[36413] = 213;
// bram[36414] = 226;
// bram[36415] = 237;
// bram[36416] = 245;
// bram[36417] = 251;
// bram[36418] = 253;
// bram[36419] = 253;
// bram[36420] = 250;
// bram[36421] = 243;
// bram[36422] = 234;
// bram[36423] = 223;
// bram[36424] = 209;
// bram[36425] = 193;
// bram[36426] = 175;
// bram[36427] = 157;
// bram[36428] = 138;
// bram[36429] = 118;
// bram[36430] = 99;
// bram[36431] = 80;
// bram[36432] = 63;
// bram[36433] = 46;
// bram[36434] = 32;
// bram[36435] = 20;
// bram[36436] = 11;
// bram[36437] = 4;
// bram[36438] = 0;
// bram[36439] = 0;
// bram[36440] = 2;
// bram[36441] = 7;
// bram[36442] = 15;
// bram[36443] = 25;
// bram[36444] = 38;
// bram[36445] = 53;
// bram[36446] = 70;
// bram[36447] = 88;
// bram[36448] = 107;
// bram[36449] = 127;
// bram[36450] = 146;
// bram[36451] = 165;
// bram[36452] = 183;
// bram[36453] = 200;
// bram[36454] = 215;
// bram[36455] = 228;
// bram[36456] = 239;
// bram[36457] = 246;
// bram[36458] = 251;
// bram[36459] = 253;
// bram[36460] = 252;
// bram[36461] = 249;
// bram[36462] = 242;
// bram[36463] = 232;
// bram[36464] = 220;
// bram[36465] = 206;
// bram[36466] = 190;
// bram[36467] = 172;
// bram[36468] = 153;
// bram[36469] = 134;
// bram[36470] = 115;
// bram[36471] = 95;
// bram[36472] = 77;
// bram[36473] = 59;
// bram[36474] = 44;
// bram[36475] = 30;
// bram[36476] = 18;
// bram[36477] = 9;
// bram[36478] = 3;
// bram[36479] = 0;
// bram[36480] = 0;
// bram[36481] = 2;
// bram[36482] = 8;
// bram[36483] = 17;
// bram[36484] = 28;
// bram[36485] = 41;
// bram[36486] = 56;
// bram[36487] = 74;
// bram[36488] = 92;
// bram[36489] = 111;
// bram[36490] = 130;
// bram[36491] = 150;
// bram[36492] = 169;
// bram[36493] = 187;
// bram[36494] = 203;
// bram[36495] = 218;
// bram[36496] = 230;
// bram[36497] = 240;
// bram[36498] = 248;
// bram[36499] = 252;
// bram[36500] = 254;
// bram[36501] = 252;
// bram[36502] = 248;
// bram[36503] = 240;
// bram[36504] = 230;
// bram[36505] = 218;
// bram[36506] = 203;
// bram[36507] = 187;
// bram[36508] = 169;
// bram[36509] = 150;
// bram[36510] = 130;
// bram[36511] = 111;
// bram[36512] = 92;
// bram[36513] = 74;
// bram[36514] = 56;
// bram[36515] = 41;
// bram[36516] = 28;
// bram[36517] = 17;
// bram[36518] = 8;
// bram[36519] = 2;
// bram[36520] = 0;
// bram[36521] = 0;
// bram[36522] = 3;
// bram[36523] = 9;
// bram[36524] = 18;
// bram[36525] = 30;
// bram[36526] = 44;
// bram[36527] = 59;
// bram[36528] = 77;
// bram[36529] = 95;
// bram[36530] = 115;
// bram[36531] = 134;
// bram[36532] = 153;
// bram[36533] = 172;
// bram[36534] = 190;
// bram[36535] = 206;
// bram[36536] = 220;
// bram[36537] = 232;
// bram[36538] = 242;
// bram[36539] = 249;
// bram[36540] = 252;
// bram[36541] = 253;
// bram[36542] = 251;
// bram[36543] = 246;
// bram[36544] = 239;
// bram[36545] = 228;
// bram[36546] = 215;
// bram[36547] = 200;
// bram[36548] = 183;
// bram[36549] = 165;
// bram[36550] = 146;
// bram[36551] = 127;
// bram[36552] = 107;
// bram[36553] = 88;
// bram[36554] = 70;
// bram[36555] = 53;
// bram[36556] = 38;
// bram[36557] = 25;
// bram[36558] = 15;
// bram[36559] = 7;
// bram[36560] = 2;
// bram[36561] = 0;
// bram[36562] = 0;
// bram[36563] = 4;
// bram[36564] = 11;
// bram[36565] = 20;
// bram[36566] = 32;
// bram[36567] = 46;
// bram[36568] = 63;
// bram[36569] = 80;
// bram[36570] = 99;
// bram[36571] = 118;
// bram[36572] = 138;
// bram[36573] = 157;
// bram[36574] = 175;
// bram[36575] = 193;
// bram[36576] = 209;
// bram[36577] = 223;
// bram[36578] = 234;
// bram[36579] = 243;
// bram[36580] = 250;
// bram[36581] = 253;
// bram[36582] = 253;
// bram[36583] = 251;
// bram[36584] = 245;
// bram[36585] = 237;
// bram[36586] = 226;
// bram[36587] = 213;
// bram[36588] = 197;
// bram[36589] = 180;
// bram[36590] = 162;
// bram[36591] = 143;
// bram[36592] = 123;
// bram[36593] = 104;
// bram[36594] = 85;
// bram[36595] = 67;
// bram[36596] = 51;
// bram[36597] = 36;
// bram[36598] = 23;
// bram[36599] = 13;
// bram[36600] = 6;
// bram[36601] = 1;
// bram[36602] = 0;
// bram[36603] = 1;
// bram[36604] = 5;
// bram[36605] = 12;
// bram[36606] = 22;
// bram[36607] = 35;
// bram[36608] = 49;
// bram[36609] = 66;
// bram[36610] = 83;
// bram[36611] = 102;
// bram[36612] = 122;
// bram[36613] = 141;
// bram[36614] = 160;
// bram[36615] = 179;
// bram[36616] = 196;
// bram[36617] = 211;
// bram[36618] = 225;
// bram[36619] = 236;
// bram[36620] = 245;
// bram[36621] = 250;
// bram[36622] = 253;
// bram[36623] = 253;
// bram[36624] = 250;
// bram[36625] = 244;
// bram[36626] = 235;
// bram[36627] = 224;
// bram[36628] = 210;
// bram[36629] = 194;
// bram[36630] = 177;
// bram[36631] = 158;
// bram[36632] = 139;
// bram[36633] = 120;
// bram[36634] = 100;
// bram[36635] = 82;
// bram[36636] = 64;
// bram[36637] = 48;
// bram[36638] = 33;
// bram[36639] = 21;
// bram[36640] = 12;
// bram[36641] = 5;
// bram[36642] = 1;
// bram[36643] = 0;
// bram[36644] = 1;
// bram[36645] = 6;
// bram[36646] = 14;
// bram[36647] = 24;
// bram[36648] = 37;
// bram[36649] = 52;
// bram[36650] = 69;
// bram[36651] = 87;
// bram[36652] = 106;
// bram[36653] = 125;
// bram[36654] = 145;
// bram[36655] = 164;
// bram[36656] = 182;
// bram[36657] = 199;
// bram[36658] = 214;
// bram[36659] = 227;
// bram[36660] = 238;
// bram[36661] = 246;
// bram[36662] = 251;
// bram[36663] = 253;
// bram[36664] = 253;
// bram[36665] = 249;
// bram[36666] = 242;
// bram[36667] = 233;
// bram[36668] = 221;
// bram[36669] = 207;
// bram[36670] = 191;
// bram[36671] = 174;
// bram[36672] = 155;
// bram[36673] = 136;
// bram[36674] = 116;
// bram[36675] = 97;
// bram[36676] = 78;
// bram[36677] = 61;
// bram[36678] = 45;
// bram[36679] = 31;
// bram[36680] = 19;
// bram[36681] = 10;
// bram[36682] = 4;
// bram[36683] = 0;
// bram[36684] = 0;
// bram[36685] = 2;
// bram[36686] = 8;
// bram[36687] = 16;
// bram[36688] = 27;
// bram[36689] = 40;
// bram[36690] = 55;
// bram[36691] = 72;
// bram[36692] = 90;
// bram[36693] = 109;
// bram[36694] = 129;
// bram[36695] = 148;
// bram[36696] = 167;
// bram[36697] = 185;
// bram[36698] = 202;
// bram[36699] = 217;
// bram[36700] = 229;
// bram[36701] = 239;
// bram[36702] = 247;
// bram[36703] = 252;
// bram[36704] = 253;
// bram[36705] = 252;
// bram[36706] = 248;
// bram[36707] = 241;
// bram[36708] = 231;
// bram[36709] = 219;
// bram[36710] = 204;
// bram[36711] = 188;
// bram[36712] = 170;
// bram[36713] = 151;
// bram[36714] = 132;
// bram[36715] = 113;
// bram[36716] = 93;
// bram[36717] = 75;
// bram[36718] = 58;
// bram[36719] = 42;
// bram[36720] = 29;
// bram[36721] = 17;
// bram[36722] = 9;
// bram[36723] = 3;
// bram[36724] = 0;
// bram[36725] = 0;
// bram[36726] = 3;
// bram[36727] = 9;
// bram[36728] = 18;
// bram[36729] = 29;
// bram[36730] = 43;
// bram[36731] = 58;
// bram[36732] = 75;
// bram[36733] = 94;
// bram[36734] = 113;
// bram[36735] = 132;
// bram[36736] = 152;
// bram[36737] = 171;
// bram[36738] = 188;
// bram[36739] = 205;
// bram[36740] = 219;
// bram[36741] = 231;
// bram[36742] = 241;
// bram[36743] = 248;
// bram[36744] = 252;
// bram[36745] = 253;
// bram[36746] = 252;
// bram[36747] = 247;
// bram[36748] = 239;
// bram[36749] = 229;
// bram[36750] = 216;
// bram[36751] = 201;
// bram[36752] = 185;
// bram[36753] = 167;
// bram[36754] = 148;
// bram[36755] = 128;
// bram[36756] = 109;
// bram[36757] = 90;
// bram[36758] = 72;
// bram[36759] = 55;
// bram[36760] = 40;
// bram[36761] = 26;
// bram[36762] = 16;
// bram[36763] = 7;
// bram[36764] = 2;
// bram[36765] = 0;
// bram[36766] = 0;
// bram[36767] = 4;
// bram[36768] = 10;
// bram[36769] = 19;
// bram[36770] = 31;
// bram[36771] = 45;
// bram[36772] = 61;
// bram[36773] = 79;
// bram[36774] = 97;
// bram[36775] = 117;
// bram[36776] = 136;
// bram[36777] = 155;
// bram[36778] = 174;
// bram[36779] = 191;
// bram[36780] = 207;
// bram[36781] = 221;
// bram[36782] = 233;
// bram[36783] = 243;
// bram[36784] = 249;
// bram[36785] = 253;
// bram[36786] = 253;
// bram[36787] = 251;
// bram[36788] = 246;
// bram[36789] = 238;
// bram[36790] = 227;
// bram[36791] = 214;
// bram[36792] = 199;
// bram[36793] = 182;
// bram[36794] = 163;
// bram[36795] = 144;
// bram[36796] = 125;
// bram[36797] = 105;
// bram[36798] = 86;
// bram[36799] = 68;
// bram[36800] = 52;
// bram[36801] = 37;
// bram[36802] = 24;
// bram[36803] = 14;
// bram[36804] = 6;
// bram[36805] = 1;
// bram[36806] = 0;
// bram[36807] = 1;
// bram[36808] = 5;
// bram[36809] = 12;
// bram[36810] = 21;
// bram[36811] = 34;
// bram[36812] = 48;
// bram[36813] = 64;
// bram[36814] = 82;
// bram[36815] = 101;
// bram[36816] = 120;
// bram[36817] = 140;
// bram[36818] = 159;
// bram[36819] = 177;
// bram[36820] = 195;
// bram[36821] = 210;
// bram[36822] = 224;
// bram[36823] = 235;
// bram[36824] = 244;
// bram[36825] = 250;
// bram[36826] = 253;
// bram[36827] = 253;
// bram[36828] = 250;
// bram[36829] = 244;
// bram[36830] = 236;
// bram[36831] = 225;
// bram[36832] = 211;
// bram[36833] = 196;
// bram[36834] = 178;
// bram[36835] = 160;
// bram[36836] = 141;
// bram[36837] = 121;
// bram[36838] = 102;
// bram[36839] = 83;
// bram[36840] = 65;
// bram[36841] = 49;
// bram[36842] = 34;
// bram[36843] = 22;
// bram[36844] = 12;
// bram[36845] = 5;
// bram[36846] = 1;
// bram[36847] = 0;
// bram[36848] = 1;
// bram[36849] = 6;
// bram[36850] = 13;
// bram[36851] = 24;
// bram[36852] = 36;
// bram[36853] = 51;
// bram[36854] = 67;
// bram[36855] = 85;
// bram[36856] = 104;
// bram[36857] = 124;
// bram[36858] = 143;
// bram[36859] = 162;
// bram[36860] = 181;
// bram[36861] = 198;
// bram[36862] = 213;
// bram[36863] = 226;
// bram[36864] = 237;
// bram[36865] = 245;
// bram[36866] = 251;
// bram[36867] = 253;
// bram[36868] = 253;
// bram[36869] = 249;
// bram[36870] = 243;
// bram[36871] = 234;
// bram[36872] = 222;
// bram[36873] = 208;
// bram[36874] = 193;
// bram[36875] = 175;
// bram[36876] = 157;
// bram[36877] = 137;
// bram[36878] = 118;
// bram[36879] = 98;
// bram[36880] = 80;
// bram[36881] = 62;
// bram[36882] = 46;
// bram[36883] = 32;
// bram[36884] = 20;
// bram[36885] = 11;
// bram[36886] = 4;
// bram[36887] = 0;
// bram[36888] = 0;
// bram[36889] = 2;
// bram[36890] = 7;
// bram[36891] = 15;
// bram[36892] = 26;
// bram[36893] = 39;
// bram[36894] = 54;
// bram[36895] = 71;
// bram[36896] = 89;
// bram[36897] = 108;
// bram[36898] = 127;
// bram[36899] = 147;
// bram[36900] = 166;
// bram[36901] = 184;
// bram[36902] = 201;
// bram[36903] = 215;
// bram[36904] = 228;
// bram[36905] = 239;
// bram[36906] = 247;
// bram[36907] = 251;
// bram[36908] = 253;
// bram[36909] = 252;
// bram[36910] = 248;
// bram[36911] = 242;
// bram[36912] = 232;
// bram[36913] = 220;
// bram[36914] = 206;
// bram[36915] = 189;
// bram[36916] = 172;
// bram[36917] = 153;
// bram[36918] = 134;
// bram[36919] = 114;
// bram[36920] = 95;
// bram[36921] = 76;
// bram[36922] = 59;
// bram[36923] = 43;
// bram[36924] = 30;
// bram[36925] = 18;
// bram[36926] = 9;
// bram[36927] = 3;
// bram[36928] = 0;
// bram[36929] = 0;
// bram[36930] = 3;
// bram[36931] = 8;
// bram[36932] = 17;
// bram[36933] = 28;
// bram[36934] = 41;
// bram[36935] = 57;
// bram[36936] = 74;
// bram[36937] = 92;
// bram[36938] = 111;
// bram[36939] = 131;
// bram[36940] = 150;
// bram[36941] = 169;
// bram[36942] = 187;
// bram[36943] = 203;
// bram[36944] = 218;
// bram[36945] = 230;
// bram[36946] = 240;
// bram[36947] = 248;
// bram[36948] = 252;
// bram[36949] = 253;
// bram[36950] = 252;
// bram[36951] = 247;
// bram[36952] = 240;
// bram[36953] = 230;
// bram[36954] = 217;
// bram[36955] = 203;
// bram[36956] = 186;
// bram[36957] = 168;
// bram[36958] = 150;
// bram[36959] = 130;
// bram[36960] = 111;
// bram[36961] = 91;
// bram[36962] = 73;
// bram[36963] = 56;
// bram[36964] = 41;
// bram[36965] = 27;
// bram[36966] = 16;
// bram[36967] = 8;
// bram[36968] = 2;
// bram[36969] = 0;
// bram[36970] = 0;
// bram[36971] = 3;
// bram[36972] = 10;
// bram[36973] = 19;
// bram[36974] = 30;
// bram[36975] = 44;
// bram[36976] = 60;
// bram[36977] = 77;
// bram[36978] = 96;
// bram[36979] = 115;
// bram[36980] = 134;
// bram[36981] = 154;
// bram[36982] = 173;
// bram[36983] = 190;
// bram[36984] = 206;
// bram[36985] = 220;
// bram[36986] = 232;
// bram[36987] = 242;
// bram[36988] = 249;
// bram[36989] = 253;
// bram[36990] = 253;
// bram[36991] = 251;
// bram[36992] = 246;
// bram[36993] = 238;
// bram[36994] = 228;
// bram[36995] = 215;
// bram[36996] = 200;
// bram[36997] = 183;
// bram[36998] = 165;
// bram[36999] = 146;
// bram[37000] = 127;
// bram[37001] = 107;
// bram[37002] = 88;
// bram[37003] = 70;
// bram[37004] = 53;
// bram[37005] = 38;
// bram[37006] = 25;
// bram[37007] = 15;
// bram[37008] = 7;
// bram[37009] = 2;
// bram[37010] = 0;
// bram[37011] = 0;
// bram[37012] = 4;
// bram[37013] = 11;
// bram[37014] = 21;
// bram[37015] = 33;
// bram[37016] = 47;
// bram[37017] = 63;
// bram[37018] = 80;
// bram[37019] = 99;
// bram[37020] = 119;
// bram[37021] = 138;
// bram[37022] = 157;
// bram[37023] = 176;
// bram[37024] = 193;
// bram[37025] = 209;
// bram[37026] = 223;
// bram[37027] = 234;
// bram[37028] = 243;
// bram[37029] = 250;
// bram[37030] = 253;
// bram[37031] = 253;
// bram[37032] = 251;
// bram[37033] = 245;
// bram[37034] = 237;
// bram[37035] = 226;
// bram[37036] = 212;
// bram[37037] = 197;
// bram[37038] = 180;
// bram[37039] = 162;
// bram[37040] = 142;
// bram[37041] = 123;
// bram[37042] = 103;
// bram[37043] = 85;
// bram[37044] = 67;
// bram[37045] = 50;
// bram[37046] = 36;
// bram[37047] = 23;
// bram[37048] = 13;
// bram[37049] = 6;
// bram[37050] = 1;
// bram[37051] = 0;
// bram[37052] = 1;
// bram[37053] = 5;
// bram[37054] = 13;
// bram[37055] = 23;
// bram[37056] = 35;
// bram[37057] = 50;
// bram[37058] = 66;
// bram[37059] = 84;
// bram[37060] = 103;
// bram[37061] = 122;
// bram[37062] = 142;
// bram[37063] = 161;
// bram[37064] = 179;
// bram[37065] = 196;
// bram[37066] = 212;
// bram[37067] = 225;
// bram[37068] = 236;
// bram[37069] = 245;
// bram[37070] = 250;
// bram[37071] = 253;
// bram[37072] = 253;
// bram[37073] = 250;
// bram[37074] = 244;
// bram[37075] = 235;
// bram[37076] = 223;
// bram[37077] = 210;
// bram[37078] = 194;
// bram[37079] = 177;
// bram[37080] = 158;
// bram[37081] = 139;
// bram[37082] = 119;
// bram[37083] = 100;
// bram[37084] = 81;
// bram[37085] = 64;
// bram[37086] = 47;
// bram[37087] = 33;
// bram[37088] = 21;
// bram[37089] = 11;
// bram[37090] = 5;
// bram[37091] = 1;
// bram[37092] = 0;
// bram[37093] = 2;
// bram[37094] = 6;
// bram[37095] = 14;
// bram[37096] = 25;
// bram[37097] = 38;
// bram[37098] = 52;
// bram[37099] = 69;
// bram[37100] = 87;
// bram[37101] = 106;
// bram[37102] = 126;
// bram[37103] = 145;
// bram[37104] = 164;
// bram[37105] = 182;
// bram[37106] = 199;
// bram[37107] = 214;
// bram[37108] = 227;
// bram[37109] = 238;
// bram[37110] = 246;
// bram[37111] = 251;
// bram[37112] = 253;
// bram[37113] = 253;
// bram[37114] = 249;
// bram[37115] = 242;
// bram[37116] = 233;
// bram[37117] = 221;
// bram[37118] = 207;
// bram[37119] = 191;
// bram[37120] = 173;
// bram[37121] = 155;
// bram[37122] = 135;
// bram[37123] = 116;
// bram[37124] = 96;
// bram[37125] = 78;
// bram[37126] = 60;
// bram[37127] = 45;
// bram[37128] = 31;
// bram[37129] = 19;
// bram[37130] = 10;
// bram[37131] = 4;
// bram[37132] = 0;
// bram[37133] = 0;
// bram[37134] = 2;
// bram[37135] = 8;
// bram[37136] = 16;
// bram[37137] = 27;
// bram[37138] = 40;
// bram[37139] = 55;
// bram[37140] = 72;
// bram[37141] = 91;
// bram[37142] = 110;
// bram[37143] = 129;
// bram[37144] = 149;
// bram[37145] = 168;
// bram[37146] = 186;
// bram[37147] = 202;
// bram[37148] = 217;
// bram[37149] = 229;
// bram[37150] = 240;
// bram[37151] = 247;
// bram[37152] = 252;
// bram[37153] = 253;
// bram[37154] = 252;
// bram[37155] = 248;
// bram[37156] = 241;
// bram[37157] = 231;
// bram[37158] = 219;
// bram[37159] = 204;
// bram[37160] = 188;
// bram[37161] = 170;
// bram[37162] = 151;
// bram[37163] = 132;
// bram[37164] = 112;
// bram[37165] = 93;
// bram[37166] = 75;
// bram[37167] = 57;
// bram[37168] = 42;
// bram[37169] = 28;
// bram[37170] = 17;
// bram[37171] = 9;
// bram[37172] = 3;
// bram[37173] = 0;
// bram[37174] = 0;
// bram[37175] = 3;
// bram[37176] = 9;
// bram[37177] = 18;
// bram[37178] = 29;
// bram[37179] = 43;
// bram[37180] = 58;
// bram[37181] = 76;
// bram[37182] = 94;
// bram[37183] = 113;
// bram[37184] = 133;
// bram[37185] = 152;
// bram[37186] = 171;
// bram[37187] = 189;
// bram[37188] = 205;
// bram[37189] = 219;
// bram[37190] = 232;
// bram[37191] = 241;
// bram[37192] = 248;
// bram[37193] = 252;
// bram[37194] = 253;
// bram[37195] = 252;
// bram[37196] = 247;
// bram[37197] = 239;
// bram[37198] = 229;
// bram[37199] = 216;
// bram[37200] = 201;
// bram[37201] = 185;
// bram[37202] = 167;
// bram[37203] = 148;
// bram[37204] = 128;
// bram[37205] = 109;
// bram[37206] = 90;
// bram[37207] = 71;
// bram[37208] = 54;
// bram[37209] = 39;
// bram[37210] = 26;
// bram[37211] = 15;
// bram[37212] = 7;
// bram[37213] = 2;
// bram[37214] = 0;
// bram[37215] = 0;
// bram[37216] = 4;
// bram[37217] = 10;
// bram[37218] = 20;
// bram[37219] = 32;
// bram[37220] = 46;
// bram[37221] = 62;
// bram[37222] = 79;
// bram[37223] = 98;
// bram[37224] = 117;
// bram[37225] = 136;
// bram[37226] = 156;
// bram[37227] = 174;
// bram[37228] = 192;
// bram[37229] = 208;
// bram[37230] = 222;
// bram[37231] = 234;
// bram[37232] = 243;
// bram[37233] = 249;
// bram[37234] = 253;
// bram[37235] = 253;
// bram[37236] = 251;
// bram[37237] = 246;
// bram[37238] = 237;
// bram[37239] = 227;
// bram[37240] = 213;
// bram[37241] = 198;
// bram[37242] = 181;
// bram[37243] = 163;
// bram[37244] = 144;
// bram[37245] = 125;
// bram[37246] = 105;
// bram[37247] = 86;
// bram[37248] = 68;
// bram[37249] = 52;
// bram[37250] = 37;
// bram[37251] = 24;
// bram[37252] = 14;
// bram[37253] = 6;
// bram[37254] = 1;
// bram[37255] = 0;
// bram[37256] = 1;
// bram[37257] = 5;
// bram[37258] = 12;
// bram[37259] = 22;
// bram[37260] = 34;
// bram[37261] = 48;
// bram[37262] = 65;
// bram[37263] = 82;
// bram[37264] = 101;
// bram[37265] = 121;
// bram[37266] = 140;
// bram[37267] = 159;
// bram[37268] = 178;
// bram[37269] = 195;
// bram[37270] = 210;
// bram[37271] = 224;
// bram[37272] = 235;
// bram[37273] = 244;
// bram[37274] = 250;
// bram[37275] = 253;
// bram[37276] = 253;
// bram[37277] = 250;
// bram[37278] = 244;
// bram[37279] = 236;
// bram[37280] = 224;
// bram[37281] = 211;
// bram[37282] = 195;
// bram[37283] = 178;
// bram[37284] = 160;
// bram[37285] = 140;
// bram[37286] = 121;
// bram[37287] = 102;
// bram[37288] = 83;
// bram[37289] = 65;
// bram[37290] = 49;
// bram[37291] = 34;
// bram[37292] = 22;
// bram[37293] = 12;
// bram[37294] = 5;
// bram[37295] = 1;
// bram[37296] = 0;
// bram[37297] = 1;
// bram[37298] = 6;
// bram[37299] = 14;
// bram[37300] = 24;
// bram[37301] = 36;
// bram[37302] = 51;
// bram[37303] = 68;
// bram[37304] = 86;
// bram[37305] = 105;
// bram[37306] = 124;
// bram[37307] = 144;
// bram[37308] = 163;
// bram[37309] = 181;
// bram[37310] = 198;
// bram[37311] = 213;
// bram[37312] = 226;
// bram[37313] = 237;
// bram[37314] = 245;
// bram[37315] = 251;
// bram[37316] = 253;
// bram[37317] = 253;
// bram[37318] = 249;
// bram[37319] = 243;
// bram[37320] = 234;
// bram[37321] = 222;
// bram[37322] = 208;
// bram[37323] = 192;
// bram[37324] = 175;
// bram[37325] = 156;
// bram[37326] = 137;
// bram[37327] = 117;
// bram[37328] = 98;
// bram[37329] = 79;
// bram[37330] = 62;
// bram[37331] = 46;
// bram[37332] = 32;
// bram[37333] = 20;
// bram[37334] = 11;
// bram[37335] = 4;
// bram[37336] = 0;
// bram[37337] = 0;
// bram[37338] = 2;
// bram[37339] = 7;
// bram[37340] = 15;
// bram[37341] = 26;
// bram[37342] = 39;
// bram[37343] = 54;
// bram[37344] = 71;
// bram[37345] = 89;
// bram[37346] = 108;
// bram[37347] = 128;
// bram[37348] = 147;
// bram[37349] = 166;
// bram[37350] = 184;
// bram[37351] = 201;
// bram[37352] = 216;
// bram[37353] = 229;
// bram[37354] = 239;
// bram[37355] = 247;
// bram[37356] = 252;
// bram[37357] = 253;
// bram[37358] = 252;
// bram[37359] = 248;
// bram[37360] = 241;
// bram[37361] = 232;
// bram[37362] = 220;
// bram[37363] = 205;
// bram[37364] = 189;
// bram[37365] = 171;
// bram[37366] = 153;
// bram[37367] = 133;
// bram[37368] = 114;
// bram[37369] = 95;
// bram[37370] = 76;
// bram[37371] = 59;
// bram[37372] = 43;
// bram[37373] = 29;
// bram[37374] = 18;
// bram[37375] = 9;
// bram[37376] = 3;
// bram[37377] = 0;
// bram[37378] = 0;
// bram[37379] = 3;
// bram[37380] = 8;
// bram[37381] = 17;
// bram[37382] = 28;
// bram[37383] = 42;
// bram[37384] = 57;
// bram[37385] = 74;
// bram[37386] = 93;
// bram[37387] = 112;
// bram[37388] = 131;
// bram[37389] = 151;
// bram[37390] = 170;
// bram[37391] = 187;
// bram[37392] = 204;
// bram[37393] = 218;
// bram[37394] = 231;
// bram[37395] = 241;
// bram[37396] = 248;
// bram[37397] = 252;
// bram[37398] = 253;
// bram[37399] = 252;
// bram[37400] = 247;
// bram[37401] = 240;
// bram[37402] = 230;
// bram[37403] = 217;
// bram[37404] = 202;
// bram[37405] = 186;
// bram[37406] = 168;
// bram[37407] = 149;
// bram[37408] = 130;
// bram[37409] = 110;
// bram[37410] = 91;
// bram[37411] = 73;
// bram[37412] = 56;
// bram[37413] = 40;
// bram[37414] = 27;
// bram[37415] = 16;
// bram[37416] = 8;
// bram[37417] = 2;
// bram[37418] = 0;
// bram[37419] = 0;
// bram[37420] = 3;
// bram[37421] = 10;
// bram[37422] = 19;
// bram[37423] = 30;
// bram[37424] = 44;
// bram[37425] = 60;
// bram[37426] = 78;
// bram[37427] = 96;
// bram[37428] = 115;
// bram[37429] = 135;
// bram[37430] = 154;
// bram[37431] = 173;
// bram[37432] = 190;
// bram[37433] = 207;
// bram[37434] = 221;
// bram[37435] = 233;
// bram[37436] = 242;
// bram[37437] = 249;
// bram[37438] = 253;
// bram[37439] = 253;
// bram[37440] = 251;
// bram[37441] = 246;
// bram[37442] = 238;
// bram[37443] = 228;
// bram[37444] = 215;
// bram[37445] = 200;
// bram[37446] = 183;
// bram[37447] = 165;
// bram[37448] = 146;
// bram[37449] = 126;
// bram[37450] = 107;
// bram[37451] = 88;
// bram[37452] = 70;
// bram[37453] = 53;
// bram[37454] = 38;
// bram[37455] = 25;
// bram[37456] = 14;
// bram[37457] = 7;
// bram[37458] = 2;
// bram[37459] = 0;
// bram[37460] = 1;
// bram[37461] = 4;
// bram[37462] = 11;
// bram[37463] = 21;
// bram[37464] = 33;
// bram[37465] = 47;
// bram[37466] = 63;
// bram[37467] = 81;
// bram[37468] = 100;
// bram[37469] = 119;
// bram[37470] = 138;
// bram[37471] = 158;
// bram[37472] = 176;
// bram[37473] = 194;
// bram[37474] = 209;
// bram[37475] = 223;
// bram[37476] = 235;
// bram[37477] = 244;
// bram[37478] = 250;
// bram[37479] = 253;
// bram[37480] = 253;
// bram[37481] = 251;
// bram[37482] = 245;
// bram[37483] = 236;
// bram[37484] = 225;
// bram[37485] = 212;
// bram[37486] = 197;
// bram[37487] = 179;
// bram[37488] = 161;
// bram[37489] = 142;
// bram[37490] = 123;
// bram[37491] = 103;
// bram[37492] = 84;
// bram[37493] = 66;
// bram[37494] = 50;
// bram[37495] = 35;
// bram[37496] = 23;
// bram[37497] = 13;
// bram[37498] = 5;
// bram[37499] = 1;
// bram[37500] = 0;
// bram[37501] = 1;
// bram[37502] = 5;
// bram[37503] = 13;
// bram[37504] = 23;
// bram[37505] = 35;
// bram[37506] = 50;
// bram[37507] = 66;
// bram[37508] = 84;
// bram[37509] = 103;
// bram[37510] = 123;
// bram[37511] = 142;
// bram[37512] = 161;
// bram[37513] = 179;
// bram[37514] = 197;
// bram[37515] = 212;
// bram[37516] = 225;
// bram[37517] = 236;
// bram[37518] = 245;
// bram[37519] = 251;
// bram[37520] = 253;
// bram[37521] = 253;
// bram[37522] = 250;
// bram[37523] = 244;
// bram[37524] = 235;
// bram[37525] = 223;
// bram[37526] = 209;
// bram[37527] = 194;
// bram[37528] = 176;
// bram[37529] = 158;
// bram[37530] = 138;
// bram[37531] = 119;
// bram[37532] = 100;
// bram[37533] = 81;
// bram[37534] = 63;
// bram[37535] = 47;
// bram[37536] = 33;
// bram[37537] = 21;
// bram[37538] = 11;
// bram[37539] = 4;
// bram[37540] = 1;
// bram[37541] = 0;
// bram[37542] = 2;
// bram[37543] = 7;
// bram[37544] = 14;
// bram[37545] = 25;
// bram[37546] = 38;
// bram[37547] = 53;
// bram[37548] = 70;
// bram[37549] = 88;
// bram[37550] = 107;
// bram[37551] = 126;
// bram[37552] = 146;
// bram[37553] = 165;
// bram[37554] = 183;
// bram[37555] = 200;
// bram[37556] = 215;
// bram[37557] = 228;
// bram[37558] = 238;
// bram[37559] = 246;
// bram[37560] = 251;
// bram[37561] = 253;
// bram[37562] = 253;
// bram[37563] = 249;
// bram[37564] = 242;
// bram[37565] = 233;
// bram[37566] = 221;
// bram[37567] = 207;
// bram[37568] = 190;
// bram[37569] = 173;
// bram[37570] = 154;
// bram[37571] = 135;
// bram[37572] = 115;
// bram[37573] = 96;
// bram[37574] = 78;
// bram[37575] = 60;
// bram[37576] = 44;
// bram[37577] = 30;
// bram[37578] = 19;
// bram[37579] = 10;
// bram[37580] = 3;
// bram[37581] = 0;
// bram[37582] = 0;
// bram[37583] = 2;
// bram[37584] = 8;
// bram[37585] = 16;
// bram[37586] = 27;
// bram[37587] = 40;
// bram[37588] = 56;
// bram[37589] = 73;
// bram[37590] = 91;
// bram[37591] = 110;
// bram[37592] = 130;
// bram[37593] = 149;
// bram[37594] = 168;
// bram[37595] = 186;
// bram[37596] = 202;
// bram[37597] = 217;
// bram[37598] = 230;
// bram[37599] = 240;
// bram[37600] = 247;
// bram[37601] = 252;
// bram[37602] = 253;
// bram[37603] = 252;
// bram[37604] = 248;
// bram[37605] = 241;
// bram[37606] = 231;
// bram[37607] = 218;
// bram[37608] = 204;
// bram[37609] = 187;
// bram[37610] = 170;
// bram[37611] = 151;
// bram[37612] = 131;
// bram[37613] = 112;
// bram[37614] = 93;
// bram[37615] = 74;
// bram[37616] = 57;
// bram[37617] = 42;
// bram[37618] = 28;
// bram[37619] = 17;
// bram[37620] = 8;
// bram[37621] = 3;
// bram[37622] = 0;
// bram[37623] = 0;
// bram[37624] = 3;
// bram[37625] = 9;
// bram[37626] = 18;
// bram[37627] = 29;
// bram[37628] = 43;
// bram[37629] = 59;
// bram[37630] = 76;
// bram[37631] = 95;
// bram[37632] = 114;
// bram[37633] = 133;
// bram[37634] = 153;
// bram[37635] = 171;
// bram[37636] = 189;
// bram[37637] = 205;
// bram[37638] = 220;
// bram[37639] = 232;
// bram[37640] = 241;
// bram[37641] = 248;
// bram[37642] = 252;
// bram[37643] = 253;
// bram[37644] = 252;
// bram[37645] = 247;
// bram[37646] = 239;
// bram[37647] = 229;
// bram[37648] = 216;
// bram[37649] = 201;
// bram[37650] = 184;
// bram[37651] = 166;
// bram[37652] = 147;
// bram[37653] = 128;
// bram[37654] = 108;
// bram[37655] = 89;
// bram[37656] = 71;
// bram[37657] = 54;
// bram[37658] = 39;
// bram[37659] = 26;
// bram[37660] = 15;
// bram[37661] = 7;
// bram[37662] = 2;
// bram[37663] = 0;
// bram[37664] = 0;
// bram[37665] = 4;
// bram[37666] = 11;
// bram[37667] = 20;
// bram[37668] = 32;
// bram[37669] = 46;
// bram[37670] = 62;
// bram[37671] = 79;
// bram[37672] = 98;
// bram[37673] = 117;
// bram[37674] = 137;
// bram[37675] = 156;
// bram[37676] = 175;
// bram[37677] = 192;
// bram[37678] = 208;
// bram[37679] = 222;
// bram[37680] = 234;
// bram[37681] = 243;
// bram[37682] = 249;
// bram[37683] = 253;
// bram[37684] = 253;
// bram[37685] = 251;
// bram[37686] = 245;
// bram[37687] = 237;
// bram[37688] = 226;
// bram[37689] = 213;
// bram[37690] = 198;
// bram[37691] = 181;
// bram[37692] = 163;
// bram[37693] = 144;
// bram[37694] = 124;
// bram[37695] = 105;
// bram[37696] = 86;
// bram[37697] = 68;
// bram[37698] = 51;
// bram[37699] = 36;
// bram[37700] = 24;
// bram[37701] = 14;
// bram[37702] = 6;
// bram[37703] = 1;
// bram[37704] = 0;
// bram[37705] = 1;
// bram[37706] = 5;
// bram[37707] = 12;
// bram[37708] = 22;
// bram[37709] = 34;
// bram[37710] = 49;
// bram[37711] = 65;
// bram[37712] = 83;
// bram[37713] = 102;
// bram[37714] = 121;
// bram[37715] = 140;
// bram[37716] = 160;
// bram[37717] = 178;
// bram[37718] = 195;
// bram[37719] = 211;
// bram[37720] = 224;
// bram[37721] = 236;
// bram[37722] = 244;
// bram[37723] = 250;
// bram[37724] = 253;
// bram[37725] = 253;
// bram[37726] = 250;
// bram[37727] = 244;
// bram[37728] = 235;
// bram[37729] = 224;
// bram[37730] = 210;
// bram[37731] = 195;
// bram[37732] = 178;
// bram[37733] = 159;
// bram[37734] = 140;
// bram[37735] = 121;
// bram[37736] = 101;
// bram[37737] = 82;
// bram[37738] = 65;
// bram[37739] = 48;
// bram[37740] = 34;
// bram[37741] = 22;
// bram[37742] = 12;
// bram[37743] = 5;
// bram[37744] = 1;
// bram[37745] = 0;
// bram[37746] = 1;
// bram[37747] = 6;
// bram[37748] = 14;
// bram[37749] = 24;
// bram[37750] = 37;
// bram[37751] = 52;
// bram[37752] = 68;
// bram[37753] = 86;
// bram[37754] = 105;
// bram[37755] = 125;
// bram[37756] = 144;
// bram[37757] = 163;
// bram[37758] = 181;
// bram[37759] = 198;
// bram[37760] = 213;
// bram[37761] = 227;
// bram[37762] = 237;
// bram[37763] = 246;
// bram[37764] = 251;
// bram[37765] = 253;
// bram[37766] = 253;
// bram[37767] = 249;
// bram[37768] = 243;
// bram[37769] = 234;
// bram[37770] = 222;
// bram[37771] = 208;
// bram[37772] = 192;
// bram[37773] = 174;
// bram[37774] = 156;
// bram[37775] = 136;
// bram[37776] = 117;
// bram[37777] = 98;
// bram[37778] = 79;
// bram[37779] = 62;
// bram[37780] = 46;
// bram[37781] = 32;
// bram[37782] = 20;
// bram[37783] = 10;
// bram[37784] = 4;
// bram[37785] = 0;
// bram[37786] = 0;
// bram[37787] = 2;
// bram[37788] = 7;
// bram[37789] = 15;
// bram[37790] = 26;
// bram[37791] = 39;
// bram[37792] = 54;
// bram[37793] = 71;
// bram[37794] = 90;
// bram[37795] = 109;
// bram[37796] = 128;
// bram[37797] = 148;
// bram[37798] = 167;
// bram[37799] = 185;
// bram[37800] = 201;
// bram[37801] = 216;
// bram[37802] = 229;
// bram[37803] = 239;
// bram[37804] = 247;
// bram[37805] = 252;
// bram[37806] = 253;
// bram[37807] = 252;
// bram[37808] = 248;
// bram[37809] = 241;
// bram[37810] = 232;
// bram[37811] = 219;
// bram[37812] = 205;
// bram[37813] = 189;
// bram[37814] = 171;
// bram[37815] = 152;
// bram[37816] = 133;
// bram[37817] = 113;
// bram[37818] = 94;
// bram[37819] = 76;
// bram[37820] = 58;
// bram[37821] = 43;
// bram[37822] = 29;
// bram[37823] = 18;
// bram[37824] = 9;
// bram[37825] = 3;
// bram[37826] = 0;
// bram[37827] = 0;
// bram[37828] = 3;
// bram[37829] = 9;
// bram[37830] = 17;
// bram[37831] = 28;
// bram[37832] = 42;
// bram[37833] = 57;
// bram[37834] = 75;
// bram[37835] = 93;
// bram[37836] = 112;
// bram[37837] = 132;
// bram[37838] = 151;
// bram[37839] = 170;
// bram[37840] = 188;
// bram[37841] = 204;
// bram[37842] = 219;
// bram[37843] = 231;
// bram[37844] = 241;
// bram[37845] = 248;
// bram[37846] = 252;
// bram[37847] = 253;
// bram[37848] = 252;
// bram[37849] = 247;
// bram[37850] = 240;
// bram[37851] = 229;
// bram[37852] = 217;
// bram[37853] = 202;
// bram[37854] = 186;
// bram[37855] = 168;
// bram[37856] = 149;
// bram[37857] = 129;
// bram[37858] = 110;
// bram[37859] = 91;
// bram[37860] = 72;
// bram[37861] = 55;
// bram[37862] = 40;
// bram[37863] = 27;
// bram[37864] = 16;
// bram[37865] = 8;
// bram[37866] = 2;
// bram[37867] = 0;
// bram[37868] = 0;
// bram[37869] = 4;
// bram[37870] = 10;
// bram[37871] = 19;
// bram[37872] = 31;
// bram[37873] = 45;
// bram[37874] = 60;
// bram[37875] = 78;
// bram[37876] = 96;
// bram[37877] = 116;
// bram[37878] = 135;
// bram[37879] = 155;
// bram[37880] = 173;
// bram[37881] = 191;
// bram[37882] = 207;
// bram[37883] = 221;
// bram[37884] = 233;
// bram[37885] = 242;
// bram[37886] = 249;
// bram[37887] = 253;
// bram[37888] = 253;
// bram[37889] = 251;
// bram[37890] = 246;
// bram[37891] = 238;
// bram[37892] = 227;
// bram[37893] = 214;
// bram[37894] = 199;
// bram[37895] = 182;
// bram[37896] = 164;
// bram[37897] = 145;
// bram[37898] = 126;
// bram[37899] = 106;
// bram[37900] = 87;
// bram[37901] = 69;
// bram[37902] = 52;
// bram[37903] = 38;
// bram[37904] = 25;
// bram[37905] = 14;
// bram[37906] = 6;
// bram[37907] = 2;
// bram[37908] = 0;
// bram[37909] = 1;
// bram[37910] = 5;
// bram[37911] = 11;
// bram[37912] = 21;
// bram[37913] = 33;
// bram[37914] = 47;
// bram[37915] = 64;
// bram[37916] = 81;
// bram[37917] = 100;
// bram[37918] = 119;
// bram[37919] = 139;
// bram[37920] = 158;
// bram[37921] = 177;
// bram[37922] = 194;
// bram[37923] = 210;
// bram[37924] = 223;
// bram[37925] = 235;
// bram[37926] = 244;
// bram[37927] = 250;
// bram[37928] = 253;
// bram[37929] = 253;
// bram[37930] = 250;
// bram[37931] = 245;
// bram[37932] = 236;
// bram[37933] = 225;
// bram[37934] = 212;
// bram[37935] = 196;
// bram[37936] = 179;
// bram[37937] = 161;
// bram[37938] = 142;
// bram[37939] = 122;
// bram[37940] = 103;
// bram[37941] = 84;
// bram[37942] = 66;
// bram[37943] = 50;
// bram[37944] = 35;
// bram[37945] = 23;
// bram[37946] = 13;
// bram[37947] = 5;
// bram[37948] = 1;
// bram[37949] = 0;
// bram[37950] = 1;
// bram[37951] = 6;
// bram[37952] = 13;
// bram[37953] = 23;
// bram[37954] = 36;
// bram[37955] = 50;
// bram[37956] = 67;
// bram[37957] = 85;
// bram[37958] = 103;
// bram[37959] = 123;
// bram[37960] = 142;
// bram[37961] = 162;
// bram[37962] = 180;
// bram[37963] = 197;
// bram[37964] = 212;
// bram[37965] = 226;
// bram[37966] = 237;
// bram[37967] = 245;
// bram[37968] = 251;
// bram[37969] = 253;
// bram[37970] = 253;
// bram[37971] = 250;
// bram[37972] = 243;
// bram[37973] = 234;
// bram[37974] = 223;
// bram[37975] = 209;
// bram[37976] = 193;
// bram[37977] = 176;
// bram[37978] = 157;
// bram[37979] = 138;
// bram[37980] = 119;
// bram[37981] = 99;
// bram[37982] = 80;
// bram[37983] = 63;
// bram[37984] = 47;
// bram[37985] = 33;
// bram[37986] = 21;
// bram[37987] = 11;
// bram[37988] = 4;
// bram[37989] = 0;
// bram[37990] = 0;
// bram[37991] = 2;
// bram[37992] = 7;
// bram[37993] = 15;
// bram[37994] = 25;
// bram[37995] = 38;
// bram[37996] = 53;
// bram[37997] = 70;
// bram[37998] = 88;
// bram[37999] = 107;
// bram[38000] = 126;
// bram[38001] = 146;
// bram[38002] = 165;
// bram[38003] = 183;
// bram[38004] = 200;
// bram[38005] = 215;
// bram[38006] = 228;
// bram[38007] = 238;
// bram[38008] = 246;
// bram[38009] = 251;
// bram[38010] = 253;
// bram[38011] = 253;
// bram[38012] = 249;
// bram[38013] = 242;
// bram[38014] = 232;
// bram[38015] = 220;
// bram[38016] = 206;
// bram[38017] = 190;
// bram[38018] = 173;
// bram[38019] = 154;
// bram[38020] = 134;
// bram[38021] = 115;
// bram[38022] = 96;
// bram[38023] = 77;
// bram[38024] = 60;
// bram[38025] = 44;
// bram[38026] = 30;
// bram[38027] = 19;
// bram[38028] = 10;
// bram[38029] = 3;
// bram[38030] = 0;
// bram[38031] = 0;
// bram[38032] = 2;
// bram[38033] = 8;
// bram[38034] = 16;
// bram[38035] = 27;
// bram[38036] = 41;
// bram[38037] = 56;
// bram[38038] = 73;
// bram[38039] = 91;
// bram[38040] = 111;
// bram[38041] = 130;
// bram[38042] = 150;
// bram[38043] = 168;
// bram[38044] = 186;
// bram[38045] = 203;
// bram[38046] = 217;
// bram[38047] = 230;
// bram[38048] = 240;
// bram[38049] = 247;
// bram[38050] = 252;
// bram[38051] = 253;
// bram[38052] = 252;
// bram[38053] = 248;
// bram[38054] = 240;
// bram[38055] = 230;
// bram[38056] = 218;
// bram[38057] = 203;
// bram[38058] = 187;
// bram[38059] = 169;
// bram[38060] = 150;
// bram[38061] = 131;
// bram[38062] = 111;
// bram[38063] = 92;
// bram[38064] = 74;
// bram[38065] = 57;
// bram[38066] = 41;
// bram[38067] = 28;
// bram[38068] = 17;
// bram[38069] = 8;
// bram[38070] = 3;
// bram[38071] = 0;
// bram[38072] = 0;
// bram[38073] = 3;
// bram[38074] = 9;
// bram[38075] = 18;
// bram[38076] = 30;
// bram[38077] = 43;
// bram[38078] = 59;
// bram[38079] = 76;
// bram[38080] = 95;
// bram[38081] = 114;
// bram[38082] = 134;
// bram[38083] = 153;
// bram[38084] = 172;
// bram[38085] = 189;
// bram[38086] = 206;
// bram[38087] = 220;
// bram[38088] = 232;
// bram[38089] = 242;
// bram[38090] = 248;
// bram[38091] = 252;
// bram[38092] = 253;
// bram[38093] = 251;
// bram[38094] = 247;
// bram[38095] = 239;
// bram[38096] = 228;
// bram[38097] = 215;
// bram[38098] = 201;
// bram[38099] = 184;
// bram[38100] = 166;
// bram[38101] = 147;
// bram[38102] = 127;
// bram[38103] = 108;
// bram[38104] = 89;
// bram[38105] = 71;
// bram[38106] = 54;
// bram[38107] = 39;
// bram[38108] = 26;
// bram[38109] = 15;
// bram[38110] = 7;
// bram[38111] = 2;
// bram[38112] = 0;
// bram[38113] = 0;
// bram[38114] = 4;
// bram[38115] = 11;
// bram[38116] = 20;
// bram[38117] = 32;
// bram[38118] = 46;
// bram[38119] = 62;
// bram[38120] = 80;
// bram[38121] = 98;
// bram[38122] = 118;
// bram[38123] = 137;
// bram[38124] = 157;
// bram[38125] = 175;
// bram[38126] = 193;
// bram[38127] = 208;
// bram[38128] = 222;
// bram[38129] = 234;
// bram[38130] = 243;
// bram[38131] = 249;
// bram[38132] = 253;
// bram[38133] = 253;
// bram[38134] = 251;
// bram[38135] = 245;
// bram[38136] = 237;
// bram[38137] = 226;
// bram[38138] = 213;
// bram[38139] = 198;
// bram[38140] = 181;
// bram[38141] = 162;
// bram[38142] = 143;
// bram[38143] = 124;
// bram[38144] = 104;
// bram[38145] = 85;
// bram[38146] = 67;
// bram[38147] = 51;
// bram[38148] = 36;
// bram[38149] = 24;
// bram[38150] = 13;
// bram[38151] = 6;
// bram[38152] = 1;
// bram[38153] = 0;
// bram[38154] = 1;
// bram[38155] = 5;
// bram[38156] = 12;
// bram[38157] = 22;
// bram[38158] = 34;
// bram[38159] = 49;
// bram[38160] = 65;
// bram[38161] = 83;
// bram[38162] = 102;
// bram[38163] = 121;
// bram[38164] = 141;
// bram[38165] = 160;
// bram[38166] = 178;
// bram[38167] = 196;
// bram[38168] = 211;
// bram[38169] = 225;
// bram[38170] = 236;
// bram[38171] = 244;
// bram[38172] = 250;
// bram[38173] = 253;
// bram[38174] = 253;
// bram[38175] = 250;
// bram[38176] = 244;
// bram[38177] = 235;
// bram[38178] = 224;
// bram[38179] = 210;
// bram[38180] = 195;
// bram[38181] = 177;
// bram[38182] = 159;
// bram[38183] = 140;
// bram[38184] = 120;
// bram[38185] = 101;
// bram[38186] = 82;
// bram[38187] = 64;
// bram[38188] = 48;
// bram[38189] = 34;
// bram[38190] = 21;
// bram[38191] = 12;
// bram[38192] = 5;
// bram[38193] = 1;
// bram[38194] = 0;
// bram[38195] = 1;
// bram[38196] = 6;
// bram[38197] = 14;
// bram[38198] = 24;
// bram[38199] = 37;
// bram[38200] = 52;
// bram[38201] = 68;
// bram[38202] = 86;
// bram[38203] = 105;
// bram[38204] = 125;
// bram[38205] = 144;
// bram[38206] = 163;
// bram[38207] = 182;
// bram[38208] = 199;
// bram[38209] = 214;
// bram[38210] = 227;
// bram[38211] = 238;
// bram[38212] = 246;
// bram[38213] = 251;
// bram[38214] = 253;
// bram[38215] = 253;
// bram[38216] = 249;
// bram[38217] = 243;
// bram[38218] = 233;
// bram[38219] = 221;
// bram[38220] = 207;
// bram[38221] = 191;
// bram[38222] = 174;
// bram[38223] = 155;
// bram[38224] = 136;
// bram[38225] = 117;
// bram[38226] = 97;
// bram[38227] = 79;
// bram[38228] = 61;
// bram[38229] = 45;
// bram[38230] = 31;
// bram[38231] = 19;
// bram[38232] = 10;
// bram[38233] = 4;
// bram[38234] = 0;
// bram[38235] = 0;
// bram[38236] = 2;
// bram[38237] = 7;
// bram[38238] = 16;
// bram[38239] = 26;
// bram[38240] = 40;
// bram[38241] = 55;
// bram[38242] = 72;
// bram[38243] = 90;
// bram[38244] = 109;
// bram[38245] = 128;
// bram[38246] = 148;
// bram[38247] = 167;
// bram[38248] = 185;
// bram[38249] = 201;
// bram[38250] = 216;
// bram[38251] = 229;
// bram[38252] = 239;
// bram[38253] = 247;
// bram[38254] = 252;
// bram[38255] = 253;
// bram[38256] = 252;
// bram[38257] = 248;
// bram[38258] = 241;
// bram[38259] = 231;
// bram[38260] = 219;
// bram[38261] = 205;
// bram[38262] = 188;
// bram[38263] = 171;
// bram[38264] = 152;
// bram[38265] = 132;
// bram[38266] = 113;
// bram[38267] = 94;
// bram[38268] = 75;
// bram[38269] = 58;
// bram[38270] = 43;
// bram[38271] = 29;
// bram[38272] = 18;
// bram[38273] = 9;
// bram[38274] = 3;
// bram[38275] = 0;
// bram[38276] = 0;
// bram[38277] = 3;
// bram[38278] = 9;
// bram[38279] = 17;
// bram[38280] = 29;
// bram[38281] = 42;
// bram[38282] = 58;
// bram[38283] = 75;
// bram[38284] = 93;
// bram[38285] = 113;
// bram[38286] = 132;
// bram[38287] = 151;
// bram[38288] = 170;
// bram[38289] = 188;
// bram[38290] = 204;
// bram[38291] = 219;
// bram[38292] = 231;
// bram[38293] = 241;
// bram[38294] = 248;
// bram[38295] = 252;
// bram[38296] = 253;
// bram[38297] = 252;
// bram[38298] = 247;
// bram[38299] = 239;
// bram[38300] = 229;
// bram[38301] = 217;
// bram[38302] = 202;
// bram[38303] = 185;
// bram[38304] = 167;
// bram[38305] = 148;
// bram[38306] = 129;
// bram[38307] = 109;
// bram[38308] = 90;
// bram[38309] = 72;
// bram[38310] = 55;
// bram[38311] = 40;
// bram[38312] = 27;
// bram[38313] = 16;
// bram[38314] = 8;
// bram[38315] = 2;
// bram[38316] = 0;
// bram[38317] = 0;
// bram[38318] = 4;
// bram[38319] = 10;
// bram[38320] = 19;
// bram[38321] = 31;
// bram[38322] = 45;
// bram[38323] = 61;
// bram[38324] = 78;
// bram[38325] = 97;
// bram[38326] = 116;
// bram[38327] = 136;
// bram[38328] = 155;
// bram[38329] = 174;
// bram[38330] = 191;
// bram[38331] = 207;
// bram[38332] = 221;
// bram[38333] = 233;
// bram[38334] = 242;
// bram[38335] = 249;
// bram[38336] = 253;
// bram[38337] = 253;
// bram[38338] = 251;
// bram[38339] = 246;
// bram[38340] = 238;
// bram[38341] = 227;
// bram[38342] = 214;
// bram[38343] = 199;
// bram[38344] = 182;
// bram[38345] = 164;
// bram[38346] = 145;
// bram[38347] = 125;
// bram[38348] = 106;
// bram[38349] = 87;
// bram[38350] = 69;
// bram[38351] = 52;
// bram[38352] = 37;
// bram[38353] = 24;
// bram[38354] = 14;
// bram[38355] = 6;
// bram[38356] = 1;
// bram[38357] = 0;
// bram[38358] = 1;
// bram[38359] = 5;
// bram[38360] = 12;
// bram[38361] = 21;
// bram[38362] = 33;
// bram[38363] = 48;
// bram[38364] = 64;
// bram[38365] = 82;
// bram[38366] = 100;
// bram[38367] = 120;
// bram[38368] = 139;
// bram[38369] = 158;
// bram[38370] = 177;
// bram[38371] = 194;
// bram[38372] = 210;
// bram[38373] = 224;
// bram[38374] = 235;
// bram[38375] = 244;
// bram[38376] = 250;
// bram[38377] = 253;
// bram[38378] = 253;
// bram[38379] = 250;
// bram[38380] = 245;
// bram[38381] = 236;
// bram[38382] = 225;
// bram[38383] = 211;
// bram[38384] = 196;
// bram[38385] = 179;
// bram[38386] = 160;
// bram[38387] = 141;
// bram[38388] = 122;
// bram[38389] = 102;
// bram[38390] = 83;
// bram[38391] = 66;
// bram[38392] = 49;
// bram[38393] = 35;
// bram[38394] = 22;
// bram[38395] = 12;
// bram[38396] = 5;
// bram[38397] = 1;
// bram[38398] = 0;
// bram[38399] = 1;
// bram[38400] = 6;
// bram[38401] = 13;
// bram[38402] = 23;
// bram[38403] = 36;
// bram[38404] = 51;
// bram[38405] = 67;
// bram[38406] = 85;
// bram[38407] = 104;
// bram[38408] = 123;
// bram[38409] = 143;
// bram[38410] = 162;
// bram[38411] = 180;
// bram[38412] = 197;
// bram[38413] = 213;
// bram[38414] = 226;
// bram[38415] = 237;
// bram[38416] = 245;
// bram[38417] = 251;
// bram[38418] = 253;
// bram[38419] = 253;
// bram[38420] = 250;
// bram[38421] = 243;
// bram[38422] = 234;
// bram[38423] = 223;
// bram[38424] = 209;
// bram[38425] = 193;
// bram[38426] = 175;
// bram[38427] = 157;
// bram[38428] = 138;
// bram[38429] = 118;
// bram[38430] = 99;
// bram[38431] = 80;
// bram[38432] = 63;
// bram[38433] = 46;
// bram[38434] = 32;
// bram[38435] = 20;
// bram[38436] = 11;
// bram[38437] = 4;
// bram[38438] = 0;
// bram[38439] = 0;
// bram[38440] = 2;
// bram[38441] = 7;
// bram[38442] = 15;
// bram[38443] = 25;
// bram[38444] = 38;
// bram[38445] = 53;
// bram[38446] = 70;
// bram[38447] = 88;
// bram[38448] = 107;
// bram[38449] = 127;
// bram[38450] = 146;
// bram[38451] = 165;
// bram[38452] = 183;
// bram[38453] = 200;
// bram[38454] = 215;
// bram[38455] = 228;
// bram[38456] = 239;
// bram[38457] = 246;
// bram[38458] = 251;
// bram[38459] = 253;
// bram[38460] = 252;
// bram[38461] = 249;
// bram[38462] = 242;
// bram[38463] = 232;
// bram[38464] = 220;
// bram[38465] = 206;
// bram[38466] = 190;
// bram[38467] = 172;
// bram[38468] = 153;
// bram[38469] = 134;
// bram[38470] = 115;
// bram[38471] = 95;
// bram[38472] = 77;
// bram[38473] = 59;
// bram[38474] = 44;
// bram[38475] = 30;
// bram[38476] = 18;
// bram[38477] = 9;
// bram[38478] = 3;
// bram[38479] = 0;
// bram[38480] = 0;
// bram[38481] = 2;
// bram[38482] = 8;
// bram[38483] = 17;
// bram[38484] = 28;
// bram[38485] = 41;
// bram[38486] = 56;
// bram[38487] = 74;
// bram[38488] = 92;
// bram[38489] = 111;
// bram[38490] = 130;
// bram[38491] = 150;
// bram[38492] = 169;
// bram[38493] = 187;
// bram[38494] = 203;
// bram[38495] = 218;
// bram[38496] = 230;
// bram[38497] = 240;
// bram[38498] = 248;
// bram[38499] = 252;
// bram[38500] = 254;
// bram[38501] = 252;
// bram[38502] = 248;
// bram[38503] = 240;
// bram[38504] = 230;
// bram[38505] = 218;
// bram[38506] = 203;
// bram[38507] = 187;
// bram[38508] = 169;
// bram[38509] = 150;
// bram[38510] = 130;
// bram[38511] = 111;
// bram[38512] = 92;
// bram[38513] = 74;
// bram[38514] = 56;
// bram[38515] = 41;
// bram[38516] = 28;
// bram[38517] = 17;
// bram[38518] = 8;
// bram[38519] = 2;
// bram[38520] = 0;
// bram[38521] = 0;
// bram[38522] = 3;
// bram[38523] = 9;
// bram[38524] = 18;
// bram[38525] = 30;
// bram[38526] = 44;
// bram[38527] = 59;
// bram[38528] = 77;
// bram[38529] = 95;
// bram[38530] = 115;
// bram[38531] = 134;
// bram[38532] = 153;
// bram[38533] = 172;
// bram[38534] = 190;
// bram[38535] = 206;
// bram[38536] = 220;
// bram[38537] = 232;
// bram[38538] = 242;
// bram[38539] = 249;
// bram[38540] = 252;
// bram[38541] = 253;
// bram[38542] = 251;
// bram[38543] = 246;
// bram[38544] = 239;
// bram[38545] = 228;
// bram[38546] = 215;
// bram[38547] = 200;
// bram[38548] = 183;
// bram[38549] = 165;
// bram[38550] = 146;
// bram[38551] = 127;
// bram[38552] = 107;
// bram[38553] = 88;
// bram[38554] = 70;
// bram[38555] = 53;
// bram[38556] = 38;
// bram[38557] = 25;
// bram[38558] = 15;
// bram[38559] = 7;
// bram[38560] = 2;
// bram[38561] = 0;
// bram[38562] = 0;
// bram[38563] = 4;
// bram[38564] = 11;
// bram[38565] = 20;
// bram[38566] = 32;
// bram[38567] = 46;
// bram[38568] = 63;
// bram[38569] = 80;
// bram[38570] = 99;
// bram[38571] = 118;
// bram[38572] = 138;
// bram[38573] = 157;
// bram[38574] = 175;
// bram[38575] = 193;
// bram[38576] = 209;
// bram[38577] = 223;
// bram[38578] = 234;
// bram[38579] = 243;
// bram[38580] = 250;
// bram[38581] = 253;
// bram[38582] = 253;
// bram[38583] = 251;
// bram[38584] = 245;
// bram[38585] = 237;
// bram[38586] = 226;
// bram[38587] = 213;
// bram[38588] = 197;
// bram[38589] = 180;
// bram[38590] = 162;
// bram[38591] = 143;
// bram[38592] = 123;
// bram[38593] = 104;
// bram[38594] = 85;
// bram[38595] = 67;
// bram[38596] = 51;
// bram[38597] = 36;
// bram[38598] = 23;
// bram[38599] = 13;
// bram[38600] = 6;
// bram[38601] = 1;
// bram[38602] = 0;
// bram[38603] = 1;
// bram[38604] = 5;
// bram[38605] = 12;
// bram[38606] = 22;
// bram[38607] = 35;
// bram[38608] = 49;
// bram[38609] = 66;
// bram[38610] = 83;
// bram[38611] = 102;
// bram[38612] = 122;
// bram[38613] = 141;
// bram[38614] = 160;
// bram[38615] = 179;
// bram[38616] = 196;
// bram[38617] = 211;
// bram[38618] = 225;
// bram[38619] = 236;
// bram[38620] = 245;
// bram[38621] = 250;
// bram[38622] = 253;
// bram[38623] = 253;
// bram[38624] = 250;
// bram[38625] = 244;
// bram[38626] = 235;
// bram[38627] = 224;
// bram[38628] = 210;
// bram[38629] = 194;
// bram[38630] = 177;
// bram[38631] = 158;
// bram[38632] = 139;
// bram[38633] = 120;
// bram[38634] = 100;
// bram[38635] = 82;
// bram[38636] = 64;
// bram[38637] = 48;
// bram[38638] = 33;
// bram[38639] = 21;
// bram[38640] = 12;
// bram[38641] = 5;
// bram[38642] = 1;
// bram[38643] = 0;
// bram[38644] = 1;
// bram[38645] = 6;
// bram[38646] = 14;
// bram[38647] = 24;
// bram[38648] = 37;
// bram[38649] = 52;
// bram[38650] = 69;
// bram[38651] = 87;
// bram[38652] = 106;
// bram[38653] = 125;
// bram[38654] = 145;
// bram[38655] = 164;
// bram[38656] = 182;
// bram[38657] = 199;
// bram[38658] = 214;
// bram[38659] = 227;
// bram[38660] = 238;
// bram[38661] = 246;
// bram[38662] = 251;
// bram[38663] = 253;
// bram[38664] = 253;
// bram[38665] = 249;
// bram[38666] = 242;
// bram[38667] = 233;
// bram[38668] = 221;
// bram[38669] = 207;
// bram[38670] = 191;
// bram[38671] = 174;
// bram[38672] = 155;
// bram[38673] = 136;
// bram[38674] = 116;
// bram[38675] = 97;
// bram[38676] = 78;
// bram[38677] = 61;
// bram[38678] = 45;
// bram[38679] = 31;
// bram[38680] = 19;
// bram[38681] = 10;
// bram[38682] = 4;
// bram[38683] = 0;
// bram[38684] = 0;
// bram[38685] = 2;
// bram[38686] = 8;
// bram[38687] = 16;
// bram[38688] = 27;
// bram[38689] = 40;
// bram[38690] = 55;
// bram[38691] = 72;
// bram[38692] = 90;
// bram[38693] = 109;
// bram[38694] = 129;
// bram[38695] = 148;
// bram[38696] = 167;
// bram[38697] = 185;
// bram[38698] = 202;
// bram[38699] = 217;
// bram[38700] = 229;
// bram[38701] = 239;
// bram[38702] = 247;
// bram[38703] = 252;
// bram[38704] = 253;
// bram[38705] = 252;
// bram[38706] = 248;
// bram[38707] = 241;
// bram[38708] = 231;
// bram[38709] = 219;
// bram[38710] = 204;
// bram[38711] = 188;
// bram[38712] = 170;
// bram[38713] = 151;
// bram[38714] = 132;
// bram[38715] = 113;
// bram[38716] = 93;
// bram[38717] = 75;
// bram[38718] = 58;
// bram[38719] = 42;
// bram[38720] = 29;
// bram[38721] = 17;
// bram[38722] = 9;
// bram[38723] = 3;
// bram[38724] = 0;
// bram[38725] = 0;
// bram[38726] = 3;
// bram[38727] = 9;
// bram[38728] = 18;
// bram[38729] = 29;
// bram[38730] = 43;
// bram[38731] = 58;
// bram[38732] = 75;
// bram[38733] = 94;
// bram[38734] = 113;
// bram[38735] = 132;
// bram[38736] = 152;
// bram[38737] = 171;
// bram[38738] = 188;
// bram[38739] = 205;
// bram[38740] = 219;
// bram[38741] = 231;
// bram[38742] = 241;
// bram[38743] = 248;
// bram[38744] = 252;
// bram[38745] = 253;
// bram[38746] = 252;
// bram[38747] = 247;
// bram[38748] = 239;
// bram[38749] = 229;
// bram[38750] = 216;
// bram[38751] = 201;
// bram[38752] = 185;
// bram[38753] = 167;
// bram[38754] = 148;
// bram[38755] = 128;
// bram[38756] = 109;
// bram[38757] = 90;
// bram[38758] = 72;
// bram[38759] = 55;
// bram[38760] = 40;
// bram[38761] = 26;
// bram[38762] = 16;
// bram[38763] = 7;
// bram[38764] = 2;
// bram[38765] = 0;
// bram[38766] = 0;
// bram[38767] = 4;
// bram[38768] = 10;
// bram[38769] = 19;
// bram[38770] = 31;
// bram[38771] = 45;
// bram[38772] = 61;
// bram[38773] = 79;
// bram[38774] = 97;
// bram[38775] = 117;
// bram[38776] = 136;
// bram[38777] = 155;
// bram[38778] = 174;
// bram[38779] = 191;
// bram[38780] = 207;
// bram[38781] = 221;
// bram[38782] = 233;
// bram[38783] = 243;
// bram[38784] = 249;
// bram[38785] = 253;
// bram[38786] = 253;
// bram[38787] = 251;
// bram[38788] = 246;
// bram[38789] = 238;
// bram[38790] = 227;
// bram[38791] = 214;
// bram[38792] = 199;
// bram[38793] = 182;
// bram[38794] = 163;
// bram[38795] = 144;
// bram[38796] = 125;
// bram[38797] = 105;
// bram[38798] = 86;
// bram[38799] = 68;
// bram[38800] = 52;
// bram[38801] = 37;
// bram[38802] = 24;
// bram[38803] = 14;
// bram[38804] = 6;
// bram[38805] = 1;
// bram[38806] = 0;
// bram[38807] = 1;
// bram[38808] = 5;
// bram[38809] = 12;
// bram[38810] = 21;
// bram[38811] = 34;
// bram[38812] = 48;
// bram[38813] = 64;
// bram[38814] = 82;
// bram[38815] = 101;
// bram[38816] = 120;
// bram[38817] = 140;
// bram[38818] = 159;
// bram[38819] = 177;
// bram[38820] = 195;
// bram[38821] = 210;
// bram[38822] = 224;
// bram[38823] = 235;
// bram[38824] = 244;
// bram[38825] = 250;
// bram[38826] = 253;
// bram[38827] = 253;
// bram[38828] = 250;
// bram[38829] = 244;
// bram[38830] = 236;
// bram[38831] = 225;
// bram[38832] = 211;
// bram[38833] = 196;
// bram[38834] = 178;
// bram[38835] = 160;
// bram[38836] = 141;
// bram[38837] = 121;
// bram[38838] = 102;
// bram[38839] = 83;
// bram[38840] = 65;
// bram[38841] = 49;
// bram[38842] = 34;
// bram[38843] = 22;
// bram[38844] = 12;
// bram[38845] = 5;
// bram[38846] = 1;
// bram[38847] = 0;
// bram[38848] = 1;
// bram[38849] = 6;
// bram[38850] = 13;
// bram[38851] = 24;
// bram[38852] = 36;
// bram[38853] = 51;
// bram[38854] = 67;
// bram[38855] = 85;
// bram[38856] = 104;
// bram[38857] = 124;
// bram[38858] = 143;
// bram[38859] = 162;
// bram[38860] = 181;
// bram[38861] = 198;
// bram[38862] = 213;
// bram[38863] = 226;
// bram[38864] = 237;
// bram[38865] = 245;
// bram[38866] = 251;
// bram[38867] = 253;
// bram[38868] = 253;
// bram[38869] = 249;
// bram[38870] = 243;
// bram[38871] = 234;
// bram[38872] = 222;
// bram[38873] = 208;
// bram[38874] = 193;
// bram[38875] = 175;
// bram[38876] = 157;
// bram[38877] = 137;
// bram[38878] = 118;
// bram[38879] = 98;
// bram[38880] = 80;
// bram[38881] = 62;
// bram[38882] = 46;
// bram[38883] = 32;
// bram[38884] = 20;
// bram[38885] = 11;
// bram[38886] = 4;
// bram[38887] = 0;
// bram[38888] = 0;
// bram[38889] = 2;
// bram[38890] = 7;
// bram[38891] = 15;
// bram[38892] = 26;
// bram[38893] = 39;
// bram[38894] = 54;
// bram[38895] = 71;
// bram[38896] = 89;
// bram[38897] = 108;
// bram[38898] = 127;
// bram[38899] = 147;
// bram[38900] = 166;
// bram[38901] = 184;
// bram[38902] = 201;
// bram[38903] = 215;
// bram[38904] = 228;
// bram[38905] = 239;
// bram[38906] = 247;
// bram[38907] = 251;
// bram[38908] = 253;
// bram[38909] = 252;
// bram[38910] = 248;
// bram[38911] = 242;
// bram[38912] = 232;
// bram[38913] = 220;
// bram[38914] = 206;
// bram[38915] = 189;
// bram[38916] = 172;
// bram[38917] = 153;
// bram[38918] = 134;
// bram[38919] = 114;
// bram[38920] = 95;
// bram[38921] = 76;
// bram[38922] = 59;
// bram[38923] = 43;
// bram[38924] = 30;
// bram[38925] = 18;
// bram[38926] = 9;
// bram[38927] = 3;
// bram[38928] = 0;
// bram[38929] = 0;
// bram[38930] = 3;
// bram[38931] = 8;
// bram[38932] = 17;
// bram[38933] = 28;
// bram[38934] = 41;
// bram[38935] = 57;
// bram[38936] = 74;
// bram[38937] = 92;
// bram[38938] = 111;
// bram[38939] = 131;
// bram[38940] = 150;
// bram[38941] = 169;
// bram[38942] = 187;
// bram[38943] = 203;
// bram[38944] = 218;
// bram[38945] = 230;
// bram[38946] = 240;
// bram[38947] = 248;
// bram[38948] = 252;
// bram[38949] = 253;
// bram[38950] = 252;
// bram[38951] = 247;
// bram[38952] = 240;
// bram[38953] = 230;
// bram[38954] = 217;
// bram[38955] = 203;
// bram[38956] = 186;
// bram[38957] = 168;
// bram[38958] = 150;
// bram[38959] = 130;
// bram[38960] = 111;
// bram[38961] = 91;
// bram[38962] = 73;
// bram[38963] = 56;
// bram[38964] = 41;
// bram[38965] = 27;
// bram[38966] = 16;
// bram[38967] = 8;
// bram[38968] = 2;
// bram[38969] = 0;
// bram[38970] = 0;
// bram[38971] = 3;
// bram[38972] = 10;
// bram[38973] = 19;
// bram[38974] = 30;
// bram[38975] = 44;
// bram[38976] = 60;
// bram[38977] = 77;
// bram[38978] = 96;
// bram[38979] = 115;
// bram[38980] = 134;
// bram[38981] = 154;
// bram[38982] = 173;
// bram[38983] = 190;
// bram[38984] = 206;
// bram[38985] = 220;
// bram[38986] = 232;
// bram[38987] = 242;
// bram[38988] = 249;
// bram[38989] = 253;
// bram[38990] = 253;
// bram[38991] = 251;
// bram[38992] = 246;
// bram[38993] = 238;
// bram[38994] = 228;
// bram[38995] = 215;
// bram[38996] = 200;
// bram[38997] = 183;
// bram[38998] = 165;
// bram[38999] = 146;
// bram[39000] = 127;
// bram[39001] = 107;
// bram[39002] = 88;
// bram[39003] = 70;
// bram[39004] = 53;
// bram[39005] = 38;
// bram[39006] = 25;
// bram[39007] = 15;
// bram[39008] = 7;
// bram[39009] = 2;
// bram[39010] = 0;
// bram[39011] = 0;
// bram[39012] = 4;
// bram[39013] = 11;
// bram[39014] = 21;
// bram[39015] = 33;
// bram[39016] = 47;
// bram[39017] = 63;
// bram[39018] = 80;
// bram[39019] = 99;
// bram[39020] = 119;
// bram[39021] = 138;
// bram[39022] = 157;
// bram[39023] = 176;
// bram[39024] = 193;
// bram[39025] = 209;
// bram[39026] = 223;
// bram[39027] = 234;
// bram[39028] = 243;
// bram[39029] = 250;
// bram[39030] = 253;
// bram[39031] = 253;
// bram[39032] = 251;
// bram[39033] = 245;
// bram[39034] = 237;
// bram[39035] = 226;
// bram[39036] = 212;
// bram[39037] = 197;
// bram[39038] = 180;
// bram[39039] = 162;
// bram[39040] = 142;
// bram[39041] = 123;
// bram[39042] = 103;
// bram[39043] = 85;
// bram[39044] = 67;
// bram[39045] = 50;
// bram[39046] = 36;
// bram[39047] = 23;
// bram[39048] = 13;
// bram[39049] = 6;
// bram[39050] = 1;
// bram[39051] = 0;
// bram[39052] = 1;
// bram[39053] = 5;
// bram[39054] = 13;
// bram[39055] = 23;
// bram[39056] = 35;
// bram[39057] = 50;
// bram[39058] = 66;
// bram[39059] = 84;
// bram[39060] = 103;
// bram[39061] = 122;
// bram[39062] = 142;
// bram[39063] = 161;
// bram[39064] = 179;
// bram[39065] = 196;
// bram[39066] = 212;
// bram[39067] = 225;
// bram[39068] = 236;
// bram[39069] = 245;
// bram[39070] = 250;
// bram[39071] = 253;
// bram[39072] = 253;
// bram[39073] = 250;
// bram[39074] = 244;
// bram[39075] = 235;
// bram[39076] = 223;
// bram[39077] = 210;
// bram[39078] = 194;
// bram[39079] = 177;
// bram[39080] = 158;
// bram[39081] = 139;
// bram[39082] = 119;
// bram[39083] = 100;
// bram[39084] = 81;
// bram[39085] = 64;
// bram[39086] = 47;
// bram[39087] = 33;
// bram[39088] = 21;
// bram[39089] = 11;
// bram[39090] = 5;
// bram[39091] = 1;
// bram[39092] = 0;
// bram[39093] = 2;
// bram[39094] = 6;
// bram[39095] = 14;
// bram[39096] = 25;
// bram[39097] = 38;
// bram[39098] = 52;
// bram[39099] = 69;
// bram[39100] = 87;
// bram[39101] = 106;
// bram[39102] = 126;
// bram[39103] = 145;
// bram[39104] = 164;
// bram[39105] = 182;
// bram[39106] = 199;
// bram[39107] = 214;
// bram[39108] = 227;
// bram[39109] = 238;
// bram[39110] = 246;
// bram[39111] = 251;
// bram[39112] = 253;
// bram[39113] = 253;
// bram[39114] = 249;
// bram[39115] = 242;
// bram[39116] = 233;
// bram[39117] = 221;
// bram[39118] = 207;
// bram[39119] = 191;
// bram[39120] = 173;
// bram[39121] = 155;
// bram[39122] = 135;
// bram[39123] = 116;
// bram[39124] = 96;
// bram[39125] = 78;
// bram[39126] = 60;
// bram[39127] = 45;
// bram[39128] = 31;
// bram[39129] = 19;
// bram[39130] = 10;
// bram[39131] = 4;
// bram[39132] = 0;
// bram[39133] = 0;
// bram[39134] = 2;
// bram[39135] = 8;
// bram[39136] = 16;
// bram[39137] = 27;
// bram[39138] = 40;
// bram[39139] = 55;
// bram[39140] = 72;
// bram[39141] = 91;
// bram[39142] = 110;
// bram[39143] = 129;
// bram[39144] = 149;
// bram[39145] = 168;
// bram[39146] = 186;
// bram[39147] = 202;
// bram[39148] = 217;
// bram[39149] = 229;
// bram[39150] = 240;
// bram[39151] = 247;
// bram[39152] = 252;
// bram[39153] = 253;
// bram[39154] = 252;
// bram[39155] = 248;
// bram[39156] = 241;
// bram[39157] = 231;
// bram[39158] = 219;
// bram[39159] = 204;
// bram[39160] = 188;
// bram[39161] = 170;
// bram[39162] = 151;
// bram[39163] = 132;
// bram[39164] = 112;
// bram[39165] = 93;
// bram[39166] = 75;
// bram[39167] = 57;
// bram[39168] = 42;
// bram[39169] = 28;
// bram[39170] = 17;
// bram[39171] = 9;
// bram[39172] = 3;
// bram[39173] = 0;
// bram[39174] = 0;
// bram[39175] = 3;
// bram[39176] = 9;
// bram[39177] = 18;
// bram[39178] = 29;
// bram[39179] = 43;
// bram[39180] = 58;
// bram[39181] = 76;
// bram[39182] = 94;
// bram[39183] = 113;
// bram[39184] = 133;
// bram[39185] = 152;
// bram[39186] = 171;
// bram[39187] = 189;
// bram[39188] = 205;
// bram[39189] = 219;
// bram[39190] = 232;
// bram[39191] = 241;
// bram[39192] = 248;
// bram[39193] = 252;
// bram[39194] = 253;
// bram[39195] = 252;
// bram[39196] = 247;
// bram[39197] = 239;
// bram[39198] = 229;
// bram[39199] = 216;
// bram[39200] = 201;
// bram[39201] = 185;
// bram[39202] = 167;
// bram[39203] = 148;
// bram[39204] = 128;
// bram[39205] = 109;
// bram[39206] = 90;
// bram[39207] = 71;
// bram[39208] = 54;
// bram[39209] = 39;
// bram[39210] = 26;
// bram[39211] = 15;
// bram[39212] = 7;
// bram[39213] = 2;
// bram[39214] = 0;
// bram[39215] = 0;
// bram[39216] = 4;
// bram[39217] = 10;
// bram[39218] = 20;
// bram[39219] = 32;
// bram[39220] = 46;
// bram[39221] = 62;
// bram[39222] = 79;
// bram[39223] = 98;
// bram[39224] = 117;
// bram[39225] = 136;
// bram[39226] = 156;
// bram[39227] = 174;
// bram[39228] = 192;
// bram[39229] = 208;
// bram[39230] = 222;
// bram[39231] = 234;
// bram[39232] = 243;
// bram[39233] = 249;
// bram[39234] = 253;
// bram[39235] = 253;
// bram[39236] = 251;
// bram[39237] = 246;
// bram[39238] = 237;
// bram[39239] = 227;
// bram[39240] = 213;
// bram[39241] = 198;
// bram[39242] = 181;
// bram[39243] = 163;
// bram[39244] = 144;
// bram[39245] = 125;
// bram[39246] = 105;
// bram[39247] = 86;
// bram[39248] = 68;
// bram[39249] = 52;
// bram[39250] = 37;
// bram[39251] = 24;
// bram[39252] = 14;
// bram[39253] = 6;
// bram[39254] = 1;
// bram[39255] = 0;
// bram[39256] = 1;
// bram[39257] = 5;
// bram[39258] = 12;
// bram[39259] = 22;
// bram[39260] = 34;
// bram[39261] = 48;
// bram[39262] = 65;
// bram[39263] = 82;
// bram[39264] = 101;
// bram[39265] = 121;
// bram[39266] = 140;
// bram[39267] = 159;
// bram[39268] = 178;
// bram[39269] = 195;
// bram[39270] = 210;
// bram[39271] = 224;
// bram[39272] = 235;
// bram[39273] = 244;
// bram[39274] = 250;
// bram[39275] = 253;
// bram[39276] = 253;
// bram[39277] = 250;
// bram[39278] = 244;
// bram[39279] = 236;
// bram[39280] = 224;
// bram[39281] = 211;
// bram[39282] = 195;
// bram[39283] = 178;
// bram[39284] = 160;
// bram[39285] = 140;
// bram[39286] = 121;
// bram[39287] = 102;
// bram[39288] = 83;
// bram[39289] = 65;
// bram[39290] = 49;
// bram[39291] = 34;
// bram[39292] = 22;
// bram[39293] = 12;
// bram[39294] = 5;
// bram[39295] = 1;
// bram[39296] = 0;
// bram[39297] = 1;
// bram[39298] = 6;
// bram[39299] = 14;
// bram[39300] = 24;
// bram[39301] = 36;
// bram[39302] = 51;
// bram[39303] = 68;
// bram[39304] = 86;
// bram[39305] = 105;
// bram[39306] = 124;
// bram[39307] = 144;
// bram[39308] = 163;
// bram[39309] = 181;
// bram[39310] = 198;
// bram[39311] = 213;
// bram[39312] = 226;
// bram[39313] = 237;
// bram[39314] = 245;
// bram[39315] = 251;
// bram[39316] = 253;
// bram[39317] = 253;
// bram[39318] = 249;
// bram[39319] = 243;
// bram[39320] = 234;
// bram[39321] = 222;
// bram[39322] = 208;
// bram[39323] = 192;
// bram[39324] = 175;
// bram[39325] = 156;
// bram[39326] = 137;
// bram[39327] = 117;
// bram[39328] = 98;
// bram[39329] = 79;
// bram[39330] = 62;
// bram[39331] = 46;
// bram[39332] = 32;
// bram[39333] = 20;
// bram[39334] = 11;
// bram[39335] = 4;
// bram[39336] = 0;
// bram[39337] = 0;
// bram[39338] = 2;
// bram[39339] = 7;
// bram[39340] = 15;
// bram[39341] = 26;
// bram[39342] = 39;
// bram[39343] = 54;
// bram[39344] = 71;
// bram[39345] = 89;
// bram[39346] = 108;
// bram[39347] = 128;
// bram[39348] = 147;
// bram[39349] = 166;
// bram[39350] = 184;
// bram[39351] = 201;
// bram[39352] = 216;
// bram[39353] = 229;
// bram[39354] = 239;
// bram[39355] = 247;
// bram[39356] = 252;
// bram[39357] = 253;
// bram[39358] = 252;
// bram[39359] = 248;
// bram[39360] = 241;
// bram[39361] = 232;
// bram[39362] = 220;
// bram[39363] = 205;
// bram[39364] = 189;
// bram[39365] = 171;
// bram[39366] = 153;
// bram[39367] = 133;
// bram[39368] = 114;
// bram[39369] = 95;
// bram[39370] = 76;
// bram[39371] = 59;
// bram[39372] = 43;
// bram[39373] = 29;
// bram[39374] = 18;
// bram[39375] = 9;
// bram[39376] = 3;
// bram[39377] = 0;
// bram[39378] = 0;
// bram[39379] = 3;
// bram[39380] = 8;
// bram[39381] = 17;
// bram[39382] = 28;
// bram[39383] = 42;
// bram[39384] = 57;
// bram[39385] = 74;
// bram[39386] = 93;
// bram[39387] = 112;
// bram[39388] = 131;
// bram[39389] = 151;
// bram[39390] = 170;
// bram[39391] = 187;
// bram[39392] = 204;
// bram[39393] = 218;
// bram[39394] = 231;
// bram[39395] = 241;
// bram[39396] = 248;
// bram[39397] = 252;
// bram[39398] = 253;
// bram[39399] = 252;
// bram[39400] = 247;
// bram[39401] = 240;
// bram[39402] = 230;
// bram[39403] = 217;
// bram[39404] = 202;
// bram[39405] = 186;
// bram[39406] = 168;
// bram[39407] = 149;
// bram[39408] = 130;
// bram[39409] = 110;
// bram[39410] = 91;
// bram[39411] = 73;
// bram[39412] = 56;
// bram[39413] = 40;
// bram[39414] = 27;
// bram[39415] = 16;
// bram[39416] = 8;
// bram[39417] = 2;
// bram[39418] = 0;
// bram[39419] = 0;
// bram[39420] = 3;
// bram[39421] = 10;
// bram[39422] = 19;
// bram[39423] = 30;
// bram[39424] = 44;
// bram[39425] = 60;
// bram[39426] = 78;
// bram[39427] = 96;
// bram[39428] = 115;
// bram[39429] = 135;
// bram[39430] = 154;
// bram[39431] = 173;
// bram[39432] = 190;
// bram[39433] = 207;
// bram[39434] = 221;
// bram[39435] = 233;
// bram[39436] = 242;
// bram[39437] = 249;
// bram[39438] = 253;
// bram[39439] = 253;
// bram[39440] = 251;
// bram[39441] = 246;
// bram[39442] = 238;
// bram[39443] = 228;
// bram[39444] = 215;
// bram[39445] = 200;
// bram[39446] = 183;
// bram[39447] = 165;
// bram[39448] = 146;
// bram[39449] = 126;
// bram[39450] = 107;
// bram[39451] = 88;
// bram[39452] = 70;
// bram[39453] = 53;
// bram[39454] = 38;
// bram[39455] = 25;
// bram[39456] = 14;
// bram[39457] = 7;
// bram[39458] = 2;
// bram[39459] = 0;
// bram[39460] = 1;
// bram[39461] = 4;
// bram[39462] = 11;
// bram[39463] = 21;
// bram[39464] = 33;
// bram[39465] = 47;
// bram[39466] = 63;
// bram[39467] = 81;
// bram[39468] = 100;
// bram[39469] = 119;
// bram[39470] = 138;
// bram[39471] = 158;
// bram[39472] = 176;
// bram[39473] = 194;
// bram[39474] = 209;
// bram[39475] = 223;
// bram[39476] = 235;
// bram[39477] = 244;
// bram[39478] = 250;
// bram[39479] = 253;
// bram[39480] = 253;
// bram[39481] = 251;
// bram[39482] = 245;
// bram[39483] = 236;
// bram[39484] = 225;
// bram[39485] = 212;
// bram[39486] = 197;
// bram[39487] = 179;
// bram[39488] = 161;
// bram[39489] = 142;
// bram[39490] = 123;
// bram[39491] = 103;
// bram[39492] = 84;
// bram[39493] = 66;
// bram[39494] = 50;
// bram[39495] = 35;
// bram[39496] = 23;
// bram[39497] = 13;
// bram[39498] = 5;
// bram[39499] = 1;
// bram[39500] = 0;
// bram[39501] = 1;
// bram[39502] = 5;
// bram[39503] = 13;
// bram[39504] = 23;
// bram[39505] = 35;
// bram[39506] = 50;
// bram[39507] = 66;
// bram[39508] = 84;
// bram[39509] = 103;
// bram[39510] = 123;
// bram[39511] = 142;
// bram[39512] = 161;
// bram[39513] = 179;
// bram[39514] = 197;
// bram[39515] = 212;
// bram[39516] = 225;
// bram[39517] = 236;
// bram[39518] = 245;
// bram[39519] = 251;
// bram[39520] = 253;
// bram[39521] = 253;
// bram[39522] = 250;
// bram[39523] = 244;
// bram[39524] = 235;
// bram[39525] = 223;
// bram[39526] = 209;
// bram[39527] = 194;
// bram[39528] = 176;
// bram[39529] = 158;
// bram[39530] = 138;
// bram[39531] = 119;
// bram[39532] = 100;
// bram[39533] = 81;
// bram[39534] = 63;
// bram[39535] = 47;
// bram[39536] = 33;
// bram[39537] = 21;
// bram[39538] = 11;
// bram[39539] = 4;
// bram[39540] = 1;
// bram[39541] = 0;
// bram[39542] = 2;
// bram[39543] = 7;
// bram[39544] = 14;
// bram[39545] = 25;
// bram[39546] = 38;
// bram[39547] = 53;
// bram[39548] = 70;
// bram[39549] = 88;
// bram[39550] = 107;
// bram[39551] = 126;
// bram[39552] = 146;
// bram[39553] = 165;
// bram[39554] = 183;
// bram[39555] = 200;
// bram[39556] = 215;
// bram[39557] = 228;
// bram[39558] = 238;
// bram[39559] = 246;
// bram[39560] = 251;
// bram[39561] = 253;
// bram[39562] = 253;
// bram[39563] = 249;
// bram[39564] = 242;
// bram[39565] = 233;
// bram[39566] = 221;
// bram[39567] = 207;
// bram[39568] = 190;
// bram[39569] = 173;
// bram[39570] = 154;
// bram[39571] = 135;
// bram[39572] = 115;
// bram[39573] = 96;
// bram[39574] = 78;
// bram[39575] = 60;
// bram[39576] = 44;
// bram[39577] = 30;
// bram[39578] = 19;
// bram[39579] = 10;
// bram[39580] = 3;
// bram[39581] = 0;
// bram[39582] = 0;
// bram[39583] = 2;
// bram[39584] = 8;
// bram[39585] = 16;
// bram[39586] = 27;
// bram[39587] = 40;
// bram[39588] = 56;
// bram[39589] = 73;
// bram[39590] = 91;
// bram[39591] = 110;
// bram[39592] = 130;
// bram[39593] = 149;
// bram[39594] = 168;
// bram[39595] = 186;
// bram[39596] = 202;
// bram[39597] = 217;
// bram[39598] = 230;
// bram[39599] = 240;
// bram[39600] = 247;
// bram[39601] = 252;
// bram[39602] = 253;
// bram[39603] = 252;
// bram[39604] = 248;
// bram[39605] = 241;
// bram[39606] = 231;
// bram[39607] = 218;
// bram[39608] = 204;
// bram[39609] = 187;
// bram[39610] = 170;
// bram[39611] = 151;
// bram[39612] = 131;
// bram[39613] = 112;
// bram[39614] = 93;
// bram[39615] = 74;
// bram[39616] = 57;
// bram[39617] = 42;
// bram[39618] = 28;
// bram[39619] = 17;
// bram[39620] = 8;
// bram[39621] = 3;
// bram[39622] = 0;
// bram[39623] = 0;
// bram[39624] = 3;
// bram[39625] = 9;
// bram[39626] = 18;
// bram[39627] = 29;
// bram[39628] = 43;
// bram[39629] = 59;
// bram[39630] = 76;
// bram[39631] = 95;
// bram[39632] = 114;
// bram[39633] = 133;
// bram[39634] = 153;
// bram[39635] = 171;
// bram[39636] = 189;
// bram[39637] = 205;
// bram[39638] = 220;
// bram[39639] = 232;
// bram[39640] = 241;
// bram[39641] = 248;
// bram[39642] = 252;
// bram[39643] = 253;
// bram[39644] = 252;
// bram[39645] = 247;
// bram[39646] = 239;
// bram[39647] = 229;
// bram[39648] = 216;
// bram[39649] = 201;
// bram[39650] = 184;
// bram[39651] = 166;
// bram[39652] = 147;
// bram[39653] = 128;
// bram[39654] = 108;
// bram[39655] = 89;
// bram[39656] = 71;
// bram[39657] = 54;
// bram[39658] = 39;
// bram[39659] = 26;
// bram[39660] = 15;
// bram[39661] = 7;
// bram[39662] = 2;
// bram[39663] = 0;
// bram[39664] = 0;
// bram[39665] = 4;
// bram[39666] = 11;
// bram[39667] = 20;
// bram[39668] = 32;
// bram[39669] = 46;
// bram[39670] = 62;
// bram[39671] = 79;
// bram[39672] = 98;
// bram[39673] = 117;
// bram[39674] = 137;
// bram[39675] = 156;
// bram[39676] = 175;
// bram[39677] = 192;
// bram[39678] = 208;
// bram[39679] = 222;
// bram[39680] = 234;
// bram[39681] = 243;
// bram[39682] = 249;
// bram[39683] = 253;
// bram[39684] = 253;
// bram[39685] = 251;
// bram[39686] = 245;
// bram[39687] = 237;
// bram[39688] = 226;
// bram[39689] = 213;
// bram[39690] = 198;
// bram[39691] = 181;
// bram[39692] = 163;
// bram[39693] = 144;
// bram[39694] = 124;
// bram[39695] = 105;
// bram[39696] = 86;
// bram[39697] = 68;
// bram[39698] = 51;
// bram[39699] = 36;
// bram[39700] = 24;
// bram[39701] = 14;
// bram[39702] = 6;
// bram[39703] = 1;
// bram[39704] = 0;
// bram[39705] = 1;
// bram[39706] = 5;
// bram[39707] = 12;
// bram[39708] = 22;
// bram[39709] = 34;
// bram[39710] = 49;
// bram[39711] = 65;
// bram[39712] = 83;
// bram[39713] = 102;
// bram[39714] = 121;
// bram[39715] = 140;
// bram[39716] = 160;
// bram[39717] = 178;
// bram[39718] = 195;
// bram[39719] = 211;
// bram[39720] = 224;
// bram[39721] = 236;
// bram[39722] = 244;
// bram[39723] = 250;
// bram[39724] = 253;
// bram[39725] = 253;
// bram[39726] = 250;
// bram[39727] = 244;
// bram[39728] = 235;
// bram[39729] = 224;
// bram[39730] = 210;
// bram[39731] = 195;
// bram[39732] = 178;
// bram[39733] = 159;
// bram[39734] = 140;
// bram[39735] = 121;
// bram[39736] = 101;
// bram[39737] = 82;
// bram[39738] = 65;
// bram[39739] = 48;
// bram[39740] = 34;
// bram[39741] = 22;
// bram[39742] = 12;
// bram[39743] = 5;
// bram[39744] = 1;
// bram[39745] = 0;
// bram[39746] = 1;
// bram[39747] = 6;
// bram[39748] = 14;
// bram[39749] = 24;
// bram[39750] = 37;
// bram[39751] = 52;
// bram[39752] = 68;
// bram[39753] = 86;
// bram[39754] = 105;
// bram[39755] = 125;
// bram[39756] = 144;
// bram[39757] = 163;
// bram[39758] = 181;
// bram[39759] = 198;
// bram[39760] = 213;
// bram[39761] = 227;
// bram[39762] = 237;
// bram[39763] = 246;
// bram[39764] = 251;
// bram[39765] = 253;
// bram[39766] = 253;
// bram[39767] = 249;
// bram[39768] = 243;
// bram[39769] = 234;
// bram[39770] = 222;
// bram[39771] = 208;
// bram[39772] = 192;
// bram[39773] = 174;
// bram[39774] = 156;
// bram[39775] = 136;
// bram[39776] = 117;
// bram[39777] = 98;
// bram[39778] = 79;
// bram[39779] = 62;
// bram[39780] = 46;
// bram[39781] = 32;
// bram[39782] = 20;
// bram[39783] = 10;
// bram[39784] = 4;
// bram[39785] = 0;
// bram[39786] = 0;
// bram[39787] = 2;
// bram[39788] = 7;
// bram[39789] = 15;
// bram[39790] = 26;
// bram[39791] = 39;
// bram[39792] = 54;
// bram[39793] = 71;
// bram[39794] = 90;
// bram[39795] = 109;
// bram[39796] = 128;
// bram[39797] = 148;
// bram[39798] = 167;
// bram[39799] = 185;
// bram[39800] = 201;
// bram[39801] = 216;
// bram[39802] = 229;
// bram[39803] = 239;
// bram[39804] = 247;
// bram[39805] = 252;
// bram[39806] = 253;
// bram[39807] = 252;
// bram[39808] = 248;
// bram[39809] = 241;
// bram[39810] = 232;
// bram[39811] = 219;
// bram[39812] = 205;
// bram[39813] = 189;
// bram[39814] = 171;
// bram[39815] = 152;
// bram[39816] = 133;
// bram[39817] = 113;
// bram[39818] = 94;
// bram[39819] = 76;
// bram[39820] = 58;
// bram[39821] = 43;
// bram[39822] = 29;
// bram[39823] = 18;
// bram[39824] = 9;
// bram[39825] = 3;
// bram[39826] = 0;
// bram[39827] = 0;
// bram[39828] = 3;
// bram[39829] = 9;
// bram[39830] = 17;
// bram[39831] = 28;
// bram[39832] = 42;
// bram[39833] = 57;
// bram[39834] = 75;
// bram[39835] = 93;
// bram[39836] = 112;
// bram[39837] = 132;
// bram[39838] = 151;
// bram[39839] = 170;
// bram[39840] = 188;
// bram[39841] = 204;
// bram[39842] = 219;
// bram[39843] = 231;
// bram[39844] = 241;
// bram[39845] = 248;
// bram[39846] = 252;
// bram[39847] = 253;
// bram[39848] = 252;
// bram[39849] = 247;
// bram[39850] = 240;
// bram[39851] = 229;
// bram[39852] = 217;
// bram[39853] = 202;
// bram[39854] = 186;
// bram[39855] = 168;
// bram[39856] = 149;
// bram[39857] = 129;
// bram[39858] = 110;
// bram[39859] = 91;
// bram[39860] = 72;
// bram[39861] = 55;
// bram[39862] = 40;
// bram[39863] = 27;
// bram[39864] = 16;
// bram[39865] = 8;
// bram[39866] = 2;
// bram[39867] = 0;
// bram[39868] = 0;
// bram[39869] = 4;
// bram[39870] = 10;
// bram[39871] = 19;
// bram[39872] = 31;
// bram[39873] = 45;
// bram[39874] = 60;
// bram[39875] = 78;
// bram[39876] = 96;
// bram[39877] = 116;
// bram[39878] = 135;
// bram[39879] = 155;
// bram[39880] = 173;
// bram[39881] = 191;
// bram[39882] = 207;
// bram[39883] = 221;
// bram[39884] = 233;
// bram[39885] = 242;
// bram[39886] = 249;
// bram[39887] = 253;
// bram[39888] = 253;
// bram[39889] = 251;
// bram[39890] = 246;
// bram[39891] = 238;
// bram[39892] = 227;
// bram[39893] = 214;
// bram[39894] = 199;
// bram[39895] = 182;
// bram[39896] = 164;
// bram[39897] = 145;
// bram[39898] = 126;
// bram[39899] = 106;
// bram[39900] = 87;
// bram[39901] = 69;
// bram[39902] = 52;
// bram[39903] = 38;
// bram[39904] = 25;
// bram[39905] = 14;
// bram[39906] = 6;
// bram[39907] = 2;
// bram[39908] = 0;
// bram[39909] = 1;
// bram[39910] = 5;
// bram[39911] = 11;
// bram[39912] = 21;
// bram[39913] = 33;
// bram[39914] = 47;
// bram[39915] = 64;
// bram[39916] = 81;
// bram[39917] = 100;
// bram[39918] = 119;
// bram[39919] = 139;
// bram[39920] = 158;
// bram[39921] = 177;
// bram[39922] = 194;
// bram[39923] = 210;
// bram[39924] = 223;
// bram[39925] = 235;
// bram[39926] = 244;
// bram[39927] = 250;
// bram[39928] = 253;
// bram[39929] = 253;
// bram[39930] = 250;
// bram[39931] = 245;
// bram[39932] = 236;
// bram[39933] = 225;
// bram[39934] = 212;
// bram[39935] = 196;
// bram[39936] = 179;
// bram[39937] = 161;
// bram[39938] = 142;
// bram[39939] = 122;
// bram[39940] = 103;
// bram[39941] = 84;
// bram[39942] = 66;
// bram[39943] = 50;
// bram[39944] = 35;
// bram[39945] = 23;
// bram[39946] = 13;
// bram[39947] = 5;
// bram[39948] = 1;
// bram[39949] = 0;
// bram[39950] = 1;
// bram[39951] = 6;
// bram[39952] = 13;
// bram[39953] = 23;
// bram[39954] = 36;
// bram[39955] = 50;
// bram[39956] = 67;
// bram[39957] = 85;
// bram[39958] = 103;
// bram[39959] = 123;
// bram[39960] = 142;
// bram[39961] = 162;
// bram[39962] = 180;
// bram[39963] = 197;
// bram[39964] = 212;
// bram[39965] = 226;
// bram[39966] = 237;
// bram[39967] = 245;
// bram[39968] = 251;
// bram[39969] = 253;
// bram[39970] = 253;
// bram[39971] = 250;
// bram[39972] = 243;
// bram[39973] = 234;
// bram[39974] = 223;
// bram[39975] = 209;
// bram[39976] = 193;
// bram[39977] = 176;
// bram[39978] = 157;
// bram[39979] = 138;
// bram[39980] = 119;
// bram[39981] = 99;
// bram[39982] = 80;
// bram[39983] = 63;
// bram[39984] = 47;
// bram[39985] = 33;
// bram[39986] = 21;
// bram[39987] = 11;
// bram[39988] = 4;
// bram[39989] = 0;
// bram[39990] = 0;
// bram[39991] = 2;
// bram[39992] = 7;
// bram[39993] = 15;
// bram[39994] = 25;
// bram[39995] = 38;
// bram[39996] = 53;
// bram[39997] = 70;
// bram[39998] = 88;
// bram[39999] = 107;
// bram[40000] = 127;
// bram[40001] = 148;
// bram[40002] = 170;
// bram[40003] = 189;
// bram[40004] = 207;
// bram[40005] = 223;
// bram[40006] = 236;
// bram[40007] = 245;
// bram[40008] = 251;
// bram[40009] = 253;
// bram[40010] = 252;
// bram[40011] = 247;
// bram[40012] = 238;
// bram[40013] = 226;
// bram[40014] = 210;
// bram[40015] = 193;
// bram[40016] = 173;
// bram[40017] = 152;
// bram[40018] = 130;
// bram[40019] = 109;
// bram[40020] = 87;
// bram[40021] = 67;
// bram[40022] = 49;
// bram[40023] = 33;
// bram[40024] = 19;
// bram[40025] = 9;
// bram[40026] = 3;
// bram[40027] = 0;
// bram[40028] = 1;
// bram[40029] = 5;
// bram[40030] = 13;
// bram[40031] = 25;
// bram[40032] = 40;
// bram[40033] = 57;
// bram[40034] = 76;
// bram[40035] = 97;
// bram[40036] = 119;
// bram[40037] = 140;
// bram[40038] = 162;
// bram[40039] = 182;
// bram[40040] = 201;
// bram[40041] = 218;
// bram[40042] = 232;
// bram[40043] = 242;
// bram[40044] = 250;
// bram[40045] = 253;
// bram[40046] = 253;
// bram[40047] = 249;
// bram[40048] = 241;
// bram[40049] = 230;
// bram[40050] = 216;
// bram[40051] = 200;
// bram[40052] = 181;
// bram[40053] = 160;
// bram[40054] = 138;
// bram[40055] = 117;
// bram[40056] = 95;
// bram[40057] = 74;
// bram[40058] = 55;
// bram[40059] = 38;
// bram[40060] = 24;
// bram[40061] = 12;
// bram[40062] = 5;
// bram[40063] = 0;
// bram[40064] = 0;
// bram[40065] = 3;
// bram[40066] = 10;
// bram[40067] = 20;
// bram[40068] = 34;
// bram[40069] = 50;
// bram[40070] = 69;
// bram[40071] = 89;
// bram[40072] = 111;
// bram[40073] = 132;
// bram[40074] = 154;
// bram[40075] = 175;
// bram[40076] = 195;
// bram[40077] = 212;
// bram[40078] = 227;
// bram[40079] = 239;
// bram[40080] = 247;
// bram[40081] = 252;
// bram[40082] = 253;
// bram[40083] = 251;
// bram[40084] = 245;
// bram[40085] = 235;
// bram[40086] = 222;
// bram[40087] = 206;
// bram[40088] = 188;
// bram[40089] = 168;
// bram[40090] = 146;
// bram[40091] = 125;
// bram[40092] = 103;
// bram[40093] = 82;
// bram[40094] = 62;
// bram[40095] = 44;
// bram[40096] = 29;
// bram[40097] = 16;
// bram[40098] = 7;
// bram[40099] = 1;
// bram[40100] = 0;
// bram[40101] = 1;
// bram[40102] = 7;
// bram[40103] = 16;
// bram[40104] = 29;
// bram[40105] = 44;
// bram[40106] = 62;
// bram[40107] = 82;
// bram[40108] = 103;
// bram[40109] = 125;
// bram[40110] = 146;
// bram[40111] = 168;
// bram[40112] = 188;
// bram[40113] = 206;
// bram[40114] = 222;
// bram[40115] = 235;
// bram[40116] = 245;
// bram[40117] = 251;
// bram[40118] = 253;
// bram[40119] = 252;
// bram[40120] = 247;
// bram[40121] = 239;
// bram[40122] = 227;
// bram[40123] = 212;
// bram[40124] = 195;
// bram[40125] = 175;
// bram[40126] = 154;
// bram[40127] = 132;
// bram[40128] = 111;
// bram[40129] = 89;
// bram[40130] = 69;
// bram[40131] = 50;
// bram[40132] = 34;
// bram[40133] = 20;
// bram[40134] = 10;
// bram[40135] = 3;
// bram[40136] = 0;
// bram[40137] = 0;
// bram[40138] = 5;
// bram[40139] = 12;
// bram[40140] = 24;
// bram[40141] = 38;
// bram[40142] = 55;
// bram[40143] = 74;
// bram[40144] = 95;
// bram[40145] = 117;
// bram[40146] = 138;
// bram[40147] = 160;
// bram[40148] = 181;
// bram[40149] = 200;
// bram[40150] = 216;
// bram[40151] = 230;
// bram[40152] = 241;
// bram[40153] = 249;
// bram[40154] = 253;
// bram[40155] = 253;
// bram[40156] = 250;
// bram[40157] = 242;
// bram[40158] = 232;
// bram[40159] = 218;
// bram[40160] = 201;
// bram[40161] = 182;
// bram[40162] = 162;
// bram[40163] = 140;
// bram[40164] = 119;
// bram[40165] = 97;
// bram[40166] = 76;
// bram[40167] = 57;
// bram[40168] = 40;
// bram[40169] = 25;
// bram[40170] = 13;
// bram[40171] = 5;
// bram[40172] = 1;
// bram[40173] = 0;
// bram[40174] = 3;
// bram[40175] = 9;
// bram[40176] = 19;
// bram[40177] = 33;
// bram[40178] = 49;
// bram[40179] = 67;
// bram[40180] = 87;
// bram[40181] = 109;
// bram[40182] = 130;
// bram[40183] = 152;
// bram[40184] = 173;
// bram[40185] = 193;
// bram[40186] = 210;
// bram[40187] = 226;
// bram[40188] = 238;
// bram[40189] = 247;
// bram[40190] = 252;
// bram[40191] = 253;
// bram[40192] = 251;
// bram[40193] = 245;
// bram[40194] = 236;
// bram[40195] = 223;
// bram[40196] = 207;
// bram[40197] = 189;
// bram[40198] = 170;
// bram[40199] = 148;
// bram[40200] = 126;
// bram[40201] = 105;
// bram[40202] = 83;
// bram[40203] = 64;
// bram[40204] = 46;
// bram[40205] = 30;
// bram[40206] = 17;
// bram[40207] = 8;
// bram[40208] = 2;
// bram[40209] = 0;
// bram[40210] = 1;
// bram[40211] = 6;
// bram[40212] = 15;
// bram[40213] = 27;
// bram[40214] = 43;
// bram[40215] = 60;
// bram[40216] = 80;
// bram[40217] = 101;
// bram[40218] = 123;
// bram[40219] = 144;
// bram[40220] = 166;
// bram[40221] = 186;
// bram[40222] = 204;
// bram[40223] = 220;
// bram[40224] = 234;
// bram[40225] = 244;
// bram[40226] = 250;
// bram[40227] = 253;
// bram[40228] = 252;
// bram[40229] = 248;
// bram[40230] = 240;
// bram[40231] = 228;
// bram[40232] = 213;
// bram[40233] = 196;
// bram[40234] = 177;
// bram[40235] = 156;
// bram[40236] = 134;
// bram[40237] = 113;
// bram[40238] = 91;
// bram[40239] = 71;
// bram[40240] = 52;
// bram[40241] = 35;
// bram[40242] = 21;
// bram[40243] = 11;
// bram[40244] = 3;
// bram[40245] = 0;
// bram[40246] = 0;
// bram[40247] = 4;
// bram[40248] = 12;
// bram[40249] = 23;
// bram[40250] = 37;
// bram[40251] = 53;
// bram[40252] = 72;
// bram[40253] = 93;
// bram[40254] = 115;
// bram[40255] = 136;
// bram[40256] = 158;
// bram[40257] = 179;
// bram[40258] = 198;
// bram[40259] = 215;
// bram[40260] = 229;
// bram[40261] = 241;
// bram[40262] = 248;
// bram[40263] = 253;
// bram[40264] = 253;
// bram[40265] = 250;
// bram[40266] = 243;
// bram[40267] = 233;
// bram[40268] = 219;
// bram[40269] = 203;
// bram[40270] = 184;
// bram[40271] = 164;
// bram[40272] = 142;
// bram[40273] = 121;
// bram[40274] = 99;
// bram[40275] = 78;
// bram[40276] = 58;
// bram[40277] = 41;
// bram[40278] = 26;
// bram[40279] = 14;
// bram[40280] = 6;
// bram[40281] = 1;
// bram[40282] = 0;
// bram[40283] = 2;
// bram[40284] = 8;
// bram[40285] = 18;
// bram[40286] = 31;
// bram[40287] = 47;
// bram[40288] = 65;
// bram[40289] = 85;
// bram[40290] = 107;
// bram[40291] = 128;
// bram[40292] = 150;
// bram[40293] = 171;
// bram[40294] = 191;
// bram[40295] = 209;
// bram[40296] = 224;
// bram[40297] = 237;
// bram[40298] = 246;
// bram[40299] = 252;
// bram[40300] = 254;
// bram[40301] = 252;
// bram[40302] = 246;
// bram[40303] = 237;
// bram[40304] = 224;
// bram[40305] = 209;
// bram[40306] = 191;
// bram[40307] = 171;
// bram[40308] = 150;
// bram[40309] = 128;
// bram[40310] = 107;
// bram[40311] = 85;
// bram[40312] = 65;
// bram[40313] = 47;
// bram[40314] = 31;
// bram[40315] = 18;
// bram[40316] = 8;
// bram[40317] = 2;
// bram[40318] = 0;
// bram[40319] = 1;
// bram[40320] = 6;
// bram[40321] = 14;
// bram[40322] = 26;
// bram[40323] = 41;
// bram[40324] = 58;
// bram[40325] = 78;
// bram[40326] = 99;
// bram[40327] = 121;
// bram[40328] = 142;
// bram[40329] = 164;
// bram[40330] = 184;
// bram[40331] = 203;
// bram[40332] = 219;
// bram[40333] = 233;
// bram[40334] = 243;
// bram[40335] = 250;
// bram[40336] = 253;
// bram[40337] = 253;
// bram[40338] = 248;
// bram[40339] = 241;
// bram[40340] = 229;
// bram[40341] = 215;
// bram[40342] = 198;
// bram[40343] = 179;
// bram[40344] = 158;
// bram[40345] = 136;
// bram[40346] = 115;
// bram[40347] = 93;
// bram[40348] = 72;
// bram[40349] = 53;
// bram[40350] = 37;
// bram[40351] = 23;
// bram[40352] = 12;
// bram[40353] = 4;
// bram[40354] = 0;
// bram[40355] = 0;
// bram[40356] = 3;
// bram[40357] = 11;
// bram[40358] = 21;
// bram[40359] = 35;
// bram[40360] = 52;
// bram[40361] = 71;
// bram[40362] = 91;
// bram[40363] = 113;
// bram[40364] = 134;
// bram[40365] = 156;
// bram[40366] = 177;
// bram[40367] = 196;
// bram[40368] = 213;
// bram[40369] = 228;
// bram[40370] = 240;
// bram[40371] = 248;
// bram[40372] = 252;
// bram[40373] = 253;
// bram[40374] = 250;
// bram[40375] = 244;
// bram[40376] = 234;
// bram[40377] = 220;
// bram[40378] = 204;
// bram[40379] = 186;
// bram[40380] = 166;
// bram[40381] = 144;
// bram[40382] = 123;
// bram[40383] = 101;
// bram[40384] = 80;
// bram[40385] = 60;
// bram[40386] = 43;
// bram[40387] = 27;
// bram[40388] = 15;
// bram[40389] = 6;
// bram[40390] = 1;
// bram[40391] = 0;
// bram[40392] = 2;
// bram[40393] = 8;
// bram[40394] = 17;
// bram[40395] = 30;
// bram[40396] = 46;
// bram[40397] = 64;
// bram[40398] = 83;
// bram[40399] = 105;
// bram[40400] = 127;
// bram[40401] = 148;
// bram[40402] = 170;
// bram[40403] = 189;
// bram[40404] = 207;
// bram[40405] = 223;
// bram[40406] = 236;
// bram[40407] = 245;
// bram[40408] = 251;
// bram[40409] = 253;
// bram[40410] = 252;
// bram[40411] = 247;
// bram[40412] = 238;
// bram[40413] = 226;
// bram[40414] = 210;
// bram[40415] = 193;
// bram[40416] = 173;
// bram[40417] = 152;
// bram[40418] = 130;
// bram[40419] = 109;
// bram[40420] = 87;
// bram[40421] = 67;
// bram[40422] = 49;
// bram[40423] = 33;
// bram[40424] = 19;
// bram[40425] = 9;
// bram[40426] = 3;
// bram[40427] = 0;
// bram[40428] = 1;
// bram[40429] = 5;
// bram[40430] = 13;
// bram[40431] = 25;
// bram[40432] = 40;
// bram[40433] = 57;
// bram[40434] = 76;
// bram[40435] = 97;
// bram[40436] = 119;
// bram[40437] = 140;
// bram[40438] = 162;
// bram[40439] = 182;
// bram[40440] = 201;
// bram[40441] = 218;
// bram[40442] = 232;
// bram[40443] = 242;
// bram[40444] = 250;
// bram[40445] = 253;
// bram[40446] = 253;
// bram[40447] = 249;
// bram[40448] = 241;
// bram[40449] = 230;
// bram[40450] = 216;
// bram[40451] = 200;
// bram[40452] = 181;
// bram[40453] = 160;
// bram[40454] = 138;
// bram[40455] = 117;
// bram[40456] = 95;
// bram[40457] = 74;
// bram[40458] = 55;
// bram[40459] = 38;
// bram[40460] = 24;
// bram[40461] = 12;
// bram[40462] = 5;
// bram[40463] = 0;
// bram[40464] = 0;
// bram[40465] = 3;
// bram[40466] = 10;
// bram[40467] = 20;
// bram[40468] = 34;
// bram[40469] = 50;
// bram[40470] = 69;
// bram[40471] = 89;
// bram[40472] = 111;
// bram[40473] = 132;
// bram[40474] = 154;
// bram[40475] = 175;
// bram[40476] = 195;
// bram[40477] = 212;
// bram[40478] = 227;
// bram[40479] = 239;
// bram[40480] = 247;
// bram[40481] = 252;
// bram[40482] = 253;
// bram[40483] = 251;
// bram[40484] = 245;
// bram[40485] = 235;
// bram[40486] = 222;
// bram[40487] = 206;
// bram[40488] = 188;
// bram[40489] = 168;
// bram[40490] = 146;
// bram[40491] = 125;
// bram[40492] = 103;
// bram[40493] = 82;
// bram[40494] = 62;
// bram[40495] = 44;
// bram[40496] = 29;
// bram[40497] = 16;
// bram[40498] = 7;
// bram[40499] = 1;
// bram[40500] = 0;
// bram[40501] = 1;
// bram[40502] = 7;
// bram[40503] = 16;
// bram[40504] = 29;
// bram[40505] = 44;
// bram[40506] = 62;
// bram[40507] = 82;
// bram[40508] = 103;
// bram[40509] = 125;
// bram[40510] = 146;
// bram[40511] = 168;
// bram[40512] = 188;
// bram[40513] = 206;
// bram[40514] = 222;
// bram[40515] = 235;
// bram[40516] = 245;
// bram[40517] = 251;
// bram[40518] = 253;
// bram[40519] = 252;
// bram[40520] = 247;
// bram[40521] = 239;
// bram[40522] = 227;
// bram[40523] = 212;
// bram[40524] = 195;
// bram[40525] = 175;
// bram[40526] = 154;
// bram[40527] = 132;
// bram[40528] = 111;
// bram[40529] = 89;
// bram[40530] = 69;
// bram[40531] = 50;
// bram[40532] = 34;
// bram[40533] = 20;
// bram[40534] = 10;
// bram[40535] = 3;
// bram[40536] = 0;
// bram[40537] = 0;
// bram[40538] = 5;
// bram[40539] = 12;
// bram[40540] = 24;
// bram[40541] = 38;
// bram[40542] = 55;
// bram[40543] = 74;
// bram[40544] = 95;
// bram[40545] = 117;
// bram[40546] = 138;
// bram[40547] = 160;
// bram[40548] = 181;
// bram[40549] = 200;
// bram[40550] = 216;
// bram[40551] = 230;
// bram[40552] = 241;
// bram[40553] = 249;
// bram[40554] = 253;
// bram[40555] = 253;
// bram[40556] = 250;
// bram[40557] = 242;
// bram[40558] = 232;
// bram[40559] = 218;
// bram[40560] = 201;
// bram[40561] = 182;
// bram[40562] = 162;
// bram[40563] = 140;
// bram[40564] = 119;
// bram[40565] = 97;
// bram[40566] = 76;
// bram[40567] = 57;
// bram[40568] = 40;
// bram[40569] = 25;
// bram[40570] = 13;
// bram[40571] = 5;
// bram[40572] = 1;
// bram[40573] = 0;
// bram[40574] = 3;
// bram[40575] = 9;
// bram[40576] = 19;
// bram[40577] = 33;
// bram[40578] = 49;
// bram[40579] = 67;
// bram[40580] = 87;
// bram[40581] = 109;
// bram[40582] = 130;
// bram[40583] = 152;
// bram[40584] = 173;
// bram[40585] = 193;
// bram[40586] = 210;
// bram[40587] = 226;
// bram[40588] = 238;
// bram[40589] = 247;
// bram[40590] = 252;
// bram[40591] = 253;
// bram[40592] = 251;
// bram[40593] = 245;
// bram[40594] = 236;
// bram[40595] = 223;
// bram[40596] = 207;
// bram[40597] = 189;
// bram[40598] = 170;
// bram[40599] = 148;
// bram[40600] = 127;
// bram[40601] = 105;
// bram[40602] = 83;
// bram[40603] = 64;
// bram[40604] = 46;
// bram[40605] = 30;
// bram[40606] = 17;
// bram[40607] = 8;
// bram[40608] = 2;
// bram[40609] = 0;
// bram[40610] = 1;
// bram[40611] = 6;
// bram[40612] = 15;
// bram[40613] = 27;
// bram[40614] = 43;
// bram[40615] = 60;
// bram[40616] = 80;
// bram[40617] = 101;
// bram[40618] = 123;
// bram[40619] = 144;
// bram[40620] = 166;
// bram[40621] = 186;
// bram[40622] = 204;
// bram[40623] = 220;
// bram[40624] = 234;
// bram[40625] = 244;
// bram[40626] = 250;
// bram[40627] = 253;
// bram[40628] = 252;
// bram[40629] = 248;
// bram[40630] = 240;
// bram[40631] = 228;
// bram[40632] = 213;
// bram[40633] = 196;
// bram[40634] = 177;
// bram[40635] = 156;
// bram[40636] = 134;
// bram[40637] = 113;
// bram[40638] = 91;
// bram[40639] = 71;
// bram[40640] = 52;
// bram[40641] = 35;
// bram[40642] = 21;
// bram[40643] = 11;
// bram[40644] = 3;
// bram[40645] = 0;
// bram[40646] = 0;
// bram[40647] = 4;
// bram[40648] = 12;
// bram[40649] = 23;
// bram[40650] = 37;
// bram[40651] = 53;
// bram[40652] = 72;
// bram[40653] = 93;
// bram[40654] = 115;
// bram[40655] = 136;
// bram[40656] = 158;
// bram[40657] = 179;
// bram[40658] = 198;
// bram[40659] = 215;
// bram[40660] = 229;
// bram[40661] = 241;
// bram[40662] = 248;
// bram[40663] = 253;
// bram[40664] = 253;
// bram[40665] = 250;
// bram[40666] = 243;
// bram[40667] = 233;
// bram[40668] = 219;
// bram[40669] = 203;
// bram[40670] = 184;
// bram[40671] = 164;
// bram[40672] = 142;
// bram[40673] = 121;
// bram[40674] = 99;
// bram[40675] = 78;
// bram[40676] = 58;
// bram[40677] = 41;
// bram[40678] = 26;
// bram[40679] = 14;
// bram[40680] = 6;
// bram[40681] = 1;
// bram[40682] = 0;
// bram[40683] = 2;
// bram[40684] = 8;
// bram[40685] = 18;
// bram[40686] = 31;
// bram[40687] = 47;
// bram[40688] = 65;
// bram[40689] = 85;
// bram[40690] = 107;
// bram[40691] = 128;
// bram[40692] = 150;
// bram[40693] = 171;
// bram[40694] = 191;
// bram[40695] = 209;
// bram[40696] = 224;
// bram[40697] = 237;
// bram[40698] = 246;
// bram[40699] = 252;
// bram[40700] = 254;
// bram[40701] = 252;
// bram[40702] = 246;
// bram[40703] = 237;
// bram[40704] = 224;
// bram[40705] = 209;
// bram[40706] = 191;
// bram[40707] = 171;
// bram[40708] = 150;
// bram[40709] = 128;
// bram[40710] = 107;
// bram[40711] = 85;
// bram[40712] = 65;
// bram[40713] = 47;
// bram[40714] = 31;
// bram[40715] = 18;
// bram[40716] = 8;
// bram[40717] = 2;
// bram[40718] = 0;
// bram[40719] = 1;
// bram[40720] = 6;
// bram[40721] = 14;
// bram[40722] = 26;
// bram[40723] = 41;
// bram[40724] = 58;
// bram[40725] = 78;
// bram[40726] = 99;
// bram[40727] = 121;
// bram[40728] = 142;
// bram[40729] = 164;
// bram[40730] = 184;
// bram[40731] = 203;
// bram[40732] = 219;
// bram[40733] = 233;
// bram[40734] = 243;
// bram[40735] = 250;
// bram[40736] = 253;
// bram[40737] = 253;
// bram[40738] = 248;
// bram[40739] = 241;
// bram[40740] = 229;
// bram[40741] = 215;
// bram[40742] = 198;
// bram[40743] = 179;
// bram[40744] = 158;
// bram[40745] = 136;
// bram[40746] = 115;
// bram[40747] = 93;
// bram[40748] = 72;
// bram[40749] = 53;
// bram[40750] = 37;
// bram[40751] = 23;
// bram[40752] = 12;
// bram[40753] = 4;
// bram[40754] = 0;
// bram[40755] = 0;
// bram[40756] = 3;
// bram[40757] = 11;
// bram[40758] = 21;
// bram[40759] = 35;
// bram[40760] = 52;
// bram[40761] = 71;
// bram[40762] = 91;
// bram[40763] = 113;
// bram[40764] = 134;
// bram[40765] = 156;
// bram[40766] = 177;
// bram[40767] = 196;
// bram[40768] = 213;
// bram[40769] = 228;
// bram[40770] = 240;
// bram[40771] = 248;
// bram[40772] = 252;
// bram[40773] = 253;
// bram[40774] = 250;
// bram[40775] = 244;
// bram[40776] = 234;
// bram[40777] = 220;
// bram[40778] = 204;
// bram[40779] = 186;
// bram[40780] = 166;
// bram[40781] = 144;
// bram[40782] = 123;
// bram[40783] = 101;
// bram[40784] = 80;
// bram[40785] = 60;
// bram[40786] = 43;
// bram[40787] = 27;
// bram[40788] = 15;
// bram[40789] = 6;
// bram[40790] = 1;
// bram[40791] = 0;
// bram[40792] = 2;
// bram[40793] = 8;
// bram[40794] = 17;
// bram[40795] = 30;
// bram[40796] = 46;
// bram[40797] = 64;
// bram[40798] = 83;
// bram[40799] = 105;
// bram[40800] = 127;
// bram[40801] = 148;
// bram[40802] = 170;
// bram[40803] = 189;
// bram[40804] = 207;
// bram[40805] = 223;
// bram[40806] = 236;
// bram[40807] = 245;
// bram[40808] = 251;
// bram[40809] = 253;
// bram[40810] = 252;
// bram[40811] = 247;
// bram[40812] = 238;
// bram[40813] = 226;
// bram[40814] = 210;
// bram[40815] = 193;
// bram[40816] = 173;
// bram[40817] = 152;
// bram[40818] = 130;
// bram[40819] = 109;
// bram[40820] = 87;
// bram[40821] = 67;
// bram[40822] = 49;
// bram[40823] = 33;
// bram[40824] = 19;
// bram[40825] = 9;
// bram[40826] = 3;
// bram[40827] = 0;
// bram[40828] = 1;
// bram[40829] = 5;
// bram[40830] = 13;
// bram[40831] = 25;
// bram[40832] = 40;
// bram[40833] = 57;
// bram[40834] = 76;
// bram[40835] = 97;
// bram[40836] = 119;
// bram[40837] = 140;
// bram[40838] = 162;
// bram[40839] = 182;
// bram[40840] = 201;
// bram[40841] = 218;
// bram[40842] = 232;
// bram[40843] = 242;
// bram[40844] = 250;
// bram[40845] = 253;
// bram[40846] = 253;
// bram[40847] = 249;
// bram[40848] = 241;
// bram[40849] = 230;
// bram[40850] = 216;
// bram[40851] = 200;
// bram[40852] = 181;
// bram[40853] = 160;
// bram[40854] = 138;
// bram[40855] = 117;
// bram[40856] = 95;
// bram[40857] = 74;
// bram[40858] = 55;
// bram[40859] = 38;
// bram[40860] = 24;
// bram[40861] = 12;
// bram[40862] = 5;
// bram[40863] = 0;
// bram[40864] = 0;
// bram[40865] = 3;
// bram[40866] = 10;
// bram[40867] = 20;
// bram[40868] = 34;
// bram[40869] = 50;
// bram[40870] = 69;
// bram[40871] = 89;
// bram[40872] = 111;
// bram[40873] = 132;
// bram[40874] = 154;
// bram[40875] = 175;
// bram[40876] = 195;
// bram[40877] = 212;
// bram[40878] = 227;
// bram[40879] = 239;
// bram[40880] = 247;
// bram[40881] = 252;
// bram[40882] = 253;
// bram[40883] = 251;
// bram[40884] = 245;
// bram[40885] = 235;
// bram[40886] = 222;
// bram[40887] = 206;
// bram[40888] = 188;
// bram[40889] = 168;
// bram[40890] = 146;
// bram[40891] = 125;
// bram[40892] = 103;
// bram[40893] = 82;
// bram[40894] = 62;
// bram[40895] = 44;
// bram[40896] = 29;
// bram[40897] = 16;
// bram[40898] = 7;
// bram[40899] = 1;
// bram[40900] = 0;
// bram[40901] = 1;
// bram[40902] = 7;
// bram[40903] = 16;
// bram[40904] = 29;
// bram[40905] = 44;
// bram[40906] = 62;
// bram[40907] = 82;
// bram[40908] = 103;
// bram[40909] = 125;
// bram[40910] = 146;
// bram[40911] = 168;
// bram[40912] = 188;
// bram[40913] = 206;
// bram[40914] = 222;
// bram[40915] = 235;
// bram[40916] = 245;
// bram[40917] = 251;
// bram[40918] = 253;
// bram[40919] = 252;
// bram[40920] = 247;
// bram[40921] = 239;
// bram[40922] = 227;
// bram[40923] = 212;
// bram[40924] = 195;
// bram[40925] = 175;
// bram[40926] = 154;
// bram[40927] = 132;
// bram[40928] = 111;
// bram[40929] = 89;
// bram[40930] = 69;
// bram[40931] = 50;
// bram[40932] = 34;
// bram[40933] = 20;
// bram[40934] = 10;
// bram[40935] = 3;
// bram[40936] = 0;
// bram[40937] = 0;
// bram[40938] = 5;
// bram[40939] = 12;
// bram[40940] = 24;
// bram[40941] = 38;
// bram[40942] = 55;
// bram[40943] = 74;
// bram[40944] = 95;
// bram[40945] = 117;
// bram[40946] = 138;
// bram[40947] = 160;
// bram[40948] = 181;
// bram[40949] = 200;
// bram[40950] = 216;
// bram[40951] = 230;
// bram[40952] = 241;
// bram[40953] = 249;
// bram[40954] = 253;
// bram[40955] = 253;
// bram[40956] = 250;
// bram[40957] = 242;
// bram[40958] = 232;
// bram[40959] = 218;
// bram[40960] = 201;
// bram[40961] = 182;
// bram[40962] = 162;
// bram[40963] = 140;
// bram[40964] = 119;
// bram[40965] = 97;
// bram[40966] = 76;
// bram[40967] = 57;
// bram[40968] = 40;
// bram[40969] = 25;
// bram[40970] = 13;
// bram[40971] = 5;
// bram[40972] = 1;
// bram[40973] = 0;
// bram[40974] = 3;
// bram[40975] = 9;
// bram[40976] = 19;
// bram[40977] = 33;
// bram[40978] = 49;
// bram[40979] = 67;
// bram[40980] = 87;
// bram[40981] = 109;
// bram[40982] = 130;
// bram[40983] = 152;
// bram[40984] = 173;
// bram[40985] = 193;
// bram[40986] = 210;
// bram[40987] = 226;
// bram[40988] = 238;
// bram[40989] = 247;
// bram[40990] = 252;
// bram[40991] = 253;
// bram[40992] = 251;
// bram[40993] = 245;
// bram[40994] = 236;
// bram[40995] = 223;
// bram[40996] = 207;
// bram[40997] = 189;
// bram[40998] = 170;
// bram[40999] = 148;
// bram[41000] = 126;
// bram[41001] = 105;
// bram[41002] = 83;
// bram[41003] = 64;
// bram[41004] = 46;
// bram[41005] = 30;
// bram[41006] = 17;
// bram[41007] = 8;
// bram[41008] = 2;
// bram[41009] = 0;
// bram[41010] = 1;
// bram[41011] = 6;
// bram[41012] = 15;
// bram[41013] = 27;
// bram[41014] = 43;
// bram[41015] = 60;
// bram[41016] = 80;
// bram[41017] = 101;
// bram[41018] = 123;
// bram[41019] = 144;
// bram[41020] = 166;
// bram[41021] = 186;
// bram[41022] = 204;
// bram[41023] = 220;
// bram[41024] = 234;
// bram[41025] = 244;
// bram[41026] = 250;
// bram[41027] = 253;
// bram[41028] = 252;
// bram[41029] = 248;
// bram[41030] = 240;
// bram[41031] = 228;
// bram[41032] = 213;
// bram[41033] = 196;
// bram[41034] = 177;
// bram[41035] = 156;
// bram[41036] = 134;
// bram[41037] = 113;
// bram[41038] = 91;
// bram[41039] = 71;
// bram[41040] = 52;
// bram[41041] = 35;
// bram[41042] = 21;
// bram[41043] = 11;
// bram[41044] = 3;
// bram[41045] = 0;
// bram[41046] = 0;
// bram[41047] = 4;
// bram[41048] = 12;
// bram[41049] = 23;
// bram[41050] = 37;
// bram[41051] = 53;
// bram[41052] = 72;
// bram[41053] = 93;
// bram[41054] = 115;
// bram[41055] = 136;
// bram[41056] = 158;
// bram[41057] = 179;
// bram[41058] = 198;
// bram[41059] = 215;
// bram[41060] = 229;
// bram[41061] = 241;
// bram[41062] = 248;
// bram[41063] = 253;
// bram[41064] = 253;
// bram[41065] = 250;
// bram[41066] = 243;
// bram[41067] = 233;
// bram[41068] = 219;
// bram[41069] = 203;
// bram[41070] = 184;
// bram[41071] = 164;
// bram[41072] = 142;
// bram[41073] = 121;
// bram[41074] = 99;
// bram[41075] = 78;
// bram[41076] = 58;
// bram[41077] = 41;
// bram[41078] = 26;
// bram[41079] = 14;
// bram[41080] = 6;
// bram[41081] = 1;
// bram[41082] = 0;
// bram[41083] = 2;
// bram[41084] = 8;
// bram[41085] = 18;
// bram[41086] = 31;
// bram[41087] = 47;
// bram[41088] = 65;
// bram[41089] = 85;
// bram[41090] = 107;
// bram[41091] = 128;
// bram[41092] = 150;
// bram[41093] = 171;
// bram[41094] = 191;
// bram[41095] = 209;
// bram[41096] = 224;
// bram[41097] = 237;
// bram[41098] = 246;
// bram[41099] = 252;
// bram[41100] = 254;
// bram[41101] = 252;
// bram[41102] = 246;
// bram[41103] = 237;
// bram[41104] = 224;
// bram[41105] = 209;
// bram[41106] = 191;
// bram[41107] = 171;
// bram[41108] = 150;
// bram[41109] = 128;
// bram[41110] = 107;
// bram[41111] = 85;
// bram[41112] = 65;
// bram[41113] = 47;
// bram[41114] = 31;
// bram[41115] = 18;
// bram[41116] = 8;
// bram[41117] = 2;
// bram[41118] = 0;
// bram[41119] = 1;
// bram[41120] = 6;
// bram[41121] = 14;
// bram[41122] = 26;
// bram[41123] = 41;
// bram[41124] = 58;
// bram[41125] = 78;
// bram[41126] = 99;
// bram[41127] = 121;
// bram[41128] = 142;
// bram[41129] = 164;
// bram[41130] = 184;
// bram[41131] = 203;
// bram[41132] = 219;
// bram[41133] = 233;
// bram[41134] = 243;
// bram[41135] = 250;
// bram[41136] = 253;
// bram[41137] = 253;
// bram[41138] = 248;
// bram[41139] = 241;
// bram[41140] = 229;
// bram[41141] = 215;
// bram[41142] = 198;
// bram[41143] = 179;
// bram[41144] = 158;
// bram[41145] = 136;
// bram[41146] = 115;
// bram[41147] = 93;
// bram[41148] = 72;
// bram[41149] = 53;
// bram[41150] = 37;
// bram[41151] = 23;
// bram[41152] = 12;
// bram[41153] = 4;
// bram[41154] = 0;
// bram[41155] = 0;
// bram[41156] = 3;
// bram[41157] = 11;
// bram[41158] = 21;
// bram[41159] = 35;
// bram[41160] = 52;
// bram[41161] = 71;
// bram[41162] = 91;
// bram[41163] = 113;
// bram[41164] = 134;
// bram[41165] = 156;
// bram[41166] = 177;
// bram[41167] = 196;
// bram[41168] = 213;
// bram[41169] = 228;
// bram[41170] = 240;
// bram[41171] = 248;
// bram[41172] = 252;
// bram[41173] = 253;
// bram[41174] = 250;
// bram[41175] = 244;
// bram[41176] = 234;
// bram[41177] = 220;
// bram[41178] = 204;
// bram[41179] = 186;
// bram[41180] = 166;
// bram[41181] = 144;
// bram[41182] = 123;
// bram[41183] = 101;
// bram[41184] = 80;
// bram[41185] = 60;
// bram[41186] = 43;
// bram[41187] = 27;
// bram[41188] = 15;
// bram[41189] = 6;
// bram[41190] = 1;
// bram[41191] = 0;
// bram[41192] = 2;
// bram[41193] = 8;
// bram[41194] = 17;
// bram[41195] = 30;
// bram[41196] = 46;
// bram[41197] = 64;
// bram[41198] = 83;
// bram[41199] = 105;
// bram[41200] = 126;
// bram[41201] = 148;
// bram[41202] = 170;
// bram[41203] = 189;
// bram[41204] = 207;
// bram[41205] = 223;
// bram[41206] = 236;
// bram[41207] = 245;
// bram[41208] = 251;
// bram[41209] = 253;
// bram[41210] = 252;
// bram[41211] = 247;
// bram[41212] = 238;
// bram[41213] = 226;
// bram[41214] = 210;
// bram[41215] = 193;
// bram[41216] = 173;
// bram[41217] = 152;
// bram[41218] = 130;
// bram[41219] = 109;
// bram[41220] = 87;
// bram[41221] = 67;
// bram[41222] = 49;
// bram[41223] = 33;
// bram[41224] = 19;
// bram[41225] = 9;
// bram[41226] = 3;
// bram[41227] = 0;
// bram[41228] = 1;
// bram[41229] = 5;
// bram[41230] = 13;
// bram[41231] = 25;
// bram[41232] = 40;
// bram[41233] = 57;
// bram[41234] = 76;
// bram[41235] = 97;
// bram[41236] = 119;
// bram[41237] = 140;
// bram[41238] = 162;
// bram[41239] = 182;
// bram[41240] = 201;
// bram[41241] = 218;
// bram[41242] = 232;
// bram[41243] = 242;
// bram[41244] = 250;
// bram[41245] = 253;
// bram[41246] = 253;
// bram[41247] = 249;
// bram[41248] = 241;
// bram[41249] = 230;
// bram[41250] = 216;
// bram[41251] = 200;
// bram[41252] = 181;
// bram[41253] = 160;
// bram[41254] = 138;
// bram[41255] = 117;
// bram[41256] = 95;
// bram[41257] = 74;
// bram[41258] = 55;
// bram[41259] = 38;
// bram[41260] = 24;
// bram[41261] = 12;
// bram[41262] = 5;
// bram[41263] = 0;
// bram[41264] = 0;
// bram[41265] = 3;
// bram[41266] = 10;
// bram[41267] = 20;
// bram[41268] = 34;
// bram[41269] = 50;
// bram[41270] = 69;
// bram[41271] = 89;
// bram[41272] = 111;
// bram[41273] = 132;
// bram[41274] = 154;
// bram[41275] = 175;
// bram[41276] = 195;
// bram[41277] = 212;
// bram[41278] = 227;
// bram[41279] = 239;
// bram[41280] = 247;
// bram[41281] = 252;
// bram[41282] = 253;
// bram[41283] = 251;
// bram[41284] = 245;
// bram[41285] = 235;
// bram[41286] = 222;
// bram[41287] = 206;
// bram[41288] = 188;
// bram[41289] = 168;
// bram[41290] = 146;
// bram[41291] = 125;
// bram[41292] = 103;
// bram[41293] = 82;
// bram[41294] = 62;
// bram[41295] = 44;
// bram[41296] = 29;
// bram[41297] = 16;
// bram[41298] = 7;
// bram[41299] = 1;
// bram[41300] = 0;
// bram[41301] = 1;
// bram[41302] = 7;
// bram[41303] = 16;
// bram[41304] = 29;
// bram[41305] = 44;
// bram[41306] = 62;
// bram[41307] = 82;
// bram[41308] = 103;
// bram[41309] = 125;
// bram[41310] = 146;
// bram[41311] = 168;
// bram[41312] = 188;
// bram[41313] = 206;
// bram[41314] = 222;
// bram[41315] = 235;
// bram[41316] = 245;
// bram[41317] = 251;
// bram[41318] = 253;
// bram[41319] = 252;
// bram[41320] = 247;
// bram[41321] = 239;
// bram[41322] = 227;
// bram[41323] = 212;
// bram[41324] = 195;
// bram[41325] = 175;
// bram[41326] = 154;
// bram[41327] = 132;
// bram[41328] = 111;
// bram[41329] = 89;
// bram[41330] = 69;
// bram[41331] = 50;
// bram[41332] = 34;
// bram[41333] = 20;
// bram[41334] = 10;
// bram[41335] = 3;
// bram[41336] = 0;
// bram[41337] = 0;
// bram[41338] = 5;
// bram[41339] = 12;
// bram[41340] = 24;
// bram[41341] = 38;
// bram[41342] = 55;
// bram[41343] = 74;
// bram[41344] = 95;
// bram[41345] = 117;
// bram[41346] = 138;
// bram[41347] = 160;
// bram[41348] = 181;
// bram[41349] = 200;
// bram[41350] = 216;
// bram[41351] = 230;
// bram[41352] = 241;
// bram[41353] = 249;
// bram[41354] = 253;
// bram[41355] = 253;
// bram[41356] = 250;
// bram[41357] = 242;
// bram[41358] = 232;
// bram[41359] = 218;
// bram[41360] = 201;
// bram[41361] = 182;
// bram[41362] = 162;
// bram[41363] = 140;
// bram[41364] = 119;
// bram[41365] = 97;
// bram[41366] = 76;
// bram[41367] = 57;
// bram[41368] = 40;
// bram[41369] = 25;
// bram[41370] = 13;
// bram[41371] = 5;
// bram[41372] = 1;
// bram[41373] = 0;
// bram[41374] = 3;
// bram[41375] = 9;
// bram[41376] = 19;
// bram[41377] = 33;
// bram[41378] = 49;
// bram[41379] = 67;
// bram[41380] = 87;
// bram[41381] = 109;
// bram[41382] = 130;
// bram[41383] = 152;
// bram[41384] = 173;
// bram[41385] = 193;
// bram[41386] = 210;
// bram[41387] = 226;
// bram[41388] = 238;
// bram[41389] = 247;
// bram[41390] = 252;
// bram[41391] = 253;
// bram[41392] = 251;
// bram[41393] = 245;
// bram[41394] = 236;
// bram[41395] = 223;
// bram[41396] = 207;
// bram[41397] = 189;
// bram[41398] = 170;
// bram[41399] = 148;
// bram[41400] = 126;
// bram[41401] = 105;
// bram[41402] = 83;
// bram[41403] = 64;
// bram[41404] = 46;
// bram[41405] = 30;
// bram[41406] = 17;
// bram[41407] = 8;
// bram[41408] = 2;
// bram[41409] = 0;
// bram[41410] = 1;
// bram[41411] = 6;
// bram[41412] = 15;
// bram[41413] = 27;
// bram[41414] = 43;
// bram[41415] = 60;
// bram[41416] = 80;
// bram[41417] = 101;
// bram[41418] = 123;
// bram[41419] = 144;
// bram[41420] = 166;
// bram[41421] = 186;
// bram[41422] = 204;
// bram[41423] = 220;
// bram[41424] = 234;
// bram[41425] = 244;
// bram[41426] = 250;
// bram[41427] = 253;
// bram[41428] = 252;
// bram[41429] = 248;
// bram[41430] = 240;
// bram[41431] = 228;
// bram[41432] = 213;
// bram[41433] = 196;
// bram[41434] = 177;
// bram[41435] = 156;
// bram[41436] = 134;
// bram[41437] = 113;
// bram[41438] = 91;
// bram[41439] = 71;
// bram[41440] = 52;
// bram[41441] = 35;
// bram[41442] = 21;
// bram[41443] = 11;
// bram[41444] = 3;
// bram[41445] = 0;
// bram[41446] = 0;
// bram[41447] = 4;
// bram[41448] = 12;
// bram[41449] = 23;
// bram[41450] = 37;
// bram[41451] = 53;
// bram[41452] = 72;
// bram[41453] = 93;
// bram[41454] = 115;
// bram[41455] = 136;
// bram[41456] = 158;
// bram[41457] = 179;
// bram[41458] = 198;
// bram[41459] = 215;
// bram[41460] = 229;
// bram[41461] = 241;
// bram[41462] = 248;
// bram[41463] = 253;
// bram[41464] = 253;
// bram[41465] = 250;
// bram[41466] = 243;
// bram[41467] = 233;
// bram[41468] = 219;
// bram[41469] = 203;
// bram[41470] = 184;
// bram[41471] = 164;
// bram[41472] = 142;
// bram[41473] = 121;
// bram[41474] = 99;
// bram[41475] = 78;
// bram[41476] = 58;
// bram[41477] = 41;
// bram[41478] = 26;
// bram[41479] = 14;
// bram[41480] = 6;
// bram[41481] = 1;
// bram[41482] = 0;
// bram[41483] = 2;
// bram[41484] = 8;
// bram[41485] = 18;
// bram[41486] = 31;
// bram[41487] = 47;
// bram[41488] = 65;
// bram[41489] = 85;
// bram[41490] = 107;
// bram[41491] = 128;
// bram[41492] = 150;
// bram[41493] = 171;
// bram[41494] = 191;
// bram[41495] = 209;
// bram[41496] = 224;
// bram[41497] = 237;
// bram[41498] = 246;
// bram[41499] = 252;
// bram[41500] = 254;
// bram[41501] = 252;
// bram[41502] = 246;
// bram[41503] = 237;
// bram[41504] = 224;
// bram[41505] = 209;
// bram[41506] = 191;
// bram[41507] = 171;
// bram[41508] = 150;
// bram[41509] = 128;
// bram[41510] = 107;
// bram[41511] = 85;
// bram[41512] = 65;
// bram[41513] = 47;
// bram[41514] = 31;
// bram[41515] = 18;
// bram[41516] = 8;
// bram[41517] = 2;
// bram[41518] = 0;
// bram[41519] = 1;
// bram[41520] = 6;
// bram[41521] = 14;
// bram[41522] = 26;
// bram[41523] = 41;
// bram[41524] = 58;
// bram[41525] = 78;
// bram[41526] = 99;
// bram[41527] = 121;
// bram[41528] = 142;
// bram[41529] = 164;
// bram[41530] = 184;
// bram[41531] = 203;
// bram[41532] = 219;
// bram[41533] = 233;
// bram[41534] = 243;
// bram[41535] = 250;
// bram[41536] = 253;
// bram[41537] = 253;
// bram[41538] = 248;
// bram[41539] = 241;
// bram[41540] = 229;
// bram[41541] = 215;
// bram[41542] = 198;
// bram[41543] = 179;
// bram[41544] = 158;
// bram[41545] = 136;
// bram[41546] = 115;
// bram[41547] = 93;
// bram[41548] = 72;
// bram[41549] = 53;
// bram[41550] = 37;
// bram[41551] = 23;
// bram[41552] = 12;
// bram[41553] = 4;
// bram[41554] = 0;
// bram[41555] = 0;
// bram[41556] = 3;
// bram[41557] = 11;
// bram[41558] = 21;
// bram[41559] = 35;
// bram[41560] = 52;
// bram[41561] = 71;
// bram[41562] = 91;
// bram[41563] = 113;
// bram[41564] = 134;
// bram[41565] = 156;
// bram[41566] = 177;
// bram[41567] = 196;
// bram[41568] = 213;
// bram[41569] = 228;
// bram[41570] = 240;
// bram[41571] = 248;
// bram[41572] = 252;
// bram[41573] = 253;
// bram[41574] = 250;
// bram[41575] = 244;
// bram[41576] = 234;
// bram[41577] = 220;
// bram[41578] = 204;
// bram[41579] = 186;
// bram[41580] = 166;
// bram[41581] = 144;
// bram[41582] = 123;
// bram[41583] = 101;
// bram[41584] = 80;
// bram[41585] = 60;
// bram[41586] = 43;
// bram[41587] = 27;
// bram[41588] = 15;
// bram[41589] = 6;
// bram[41590] = 1;
// bram[41591] = 0;
// bram[41592] = 2;
// bram[41593] = 8;
// bram[41594] = 17;
// bram[41595] = 30;
// bram[41596] = 46;
// bram[41597] = 64;
// bram[41598] = 83;
// bram[41599] = 105;
// bram[41600] = 127;
// bram[41601] = 148;
// bram[41602] = 170;
// bram[41603] = 189;
// bram[41604] = 207;
// bram[41605] = 223;
// bram[41606] = 236;
// bram[41607] = 245;
// bram[41608] = 251;
// bram[41609] = 253;
// bram[41610] = 252;
// bram[41611] = 247;
// bram[41612] = 238;
// bram[41613] = 226;
// bram[41614] = 210;
// bram[41615] = 193;
// bram[41616] = 173;
// bram[41617] = 152;
// bram[41618] = 130;
// bram[41619] = 109;
// bram[41620] = 87;
// bram[41621] = 67;
// bram[41622] = 49;
// bram[41623] = 33;
// bram[41624] = 19;
// bram[41625] = 9;
// bram[41626] = 3;
// bram[41627] = 0;
// bram[41628] = 1;
// bram[41629] = 5;
// bram[41630] = 13;
// bram[41631] = 25;
// bram[41632] = 40;
// bram[41633] = 57;
// bram[41634] = 76;
// bram[41635] = 97;
// bram[41636] = 119;
// bram[41637] = 140;
// bram[41638] = 162;
// bram[41639] = 182;
// bram[41640] = 201;
// bram[41641] = 218;
// bram[41642] = 232;
// bram[41643] = 242;
// bram[41644] = 250;
// bram[41645] = 253;
// bram[41646] = 253;
// bram[41647] = 249;
// bram[41648] = 241;
// bram[41649] = 230;
// bram[41650] = 216;
// bram[41651] = 200;
// bram[41652] = 181;
// bram[41653] = 160;
// bram[41654] = 138;
// bram[41655] = 117;
// bram[41656] = 95;
// bram[41657] = 74;
// bram[41658] = 55;
// bram[41659] = 38;
// bram[41660] = 24;
// bram[41661] = 12;
// bram[41662] = 5;
// bram[41663] = 0;
// bram[41664] = 0;
// bram[41665] = 3;
// bram[41666] = 10;
// bram[41667] = 20;
// bram[41668] = 34;
// bram[41669] = 50;
// bram[41670] = 69;
// bram[41671] = 89;
// bram[41672] = 111;
// bram[41673] = 132;
// bram[41674] = 154;
// bram[41675] = 175;
// bram[41676] = 195;
// bram[41677] = 212;
// bram[41678] = 227;
// bram[41679] = 239;
// bram[41680] = 247;
// bram[41681] = 252;
// bram[41682] = 253;
// bram[41683] = 251;
// bram[41684] = 245;
// bram[41685] = 235;
// bram[41686] = 222;
// bram[41687] = 206;
// bram[41688] = 188;
// bram[41689] = 168;
// bram[41690] = 146;
// bram[41691] = 125;
// bram[41692] = 103;
// bram[41693] = 82;
// bram[41694] = 62;
// bram[41695] = 44;
// bram[41696] = 29;
// bram[41697] = 16;
// bram[41698] = 7;
// bram[41699] = 1;
// bram[41700] = 0;
// bram[41701] = 1;
// bram[41702] = 7;
// bram[41703] = 16;
// bram[41704] = 29;
// bram[41705] = 44;
// bram[41706] = 62;
// bram[41707] = 82;
// bram[41708] = 103;
// bram[41709] = 125;
// bram[41710] = 146;
// bram[41711] = 168;
// bram[41712] = 188;
// bram[41713] = 206;
// bram[41714] = 222;
// bram[41715] = 235;
// bram[41716] = 245;
// bram[41717] = 251;
// bram[41718] = 253;
// bram[41719] = 252;
// bram[41720] = 247;
// bram[41721] = 239;
// bram[41722] = 227;
// bram[41723] = 212;
// bram[41724] = 195;
// bram[41725] = 175;
// bram[41726] = 154;
// bram[41727] = 132;
// bram[41728] = 111;
// bram[41729] = 89;
// bram[41730] = 69;
// bram[41731] = 50;
// bram[41732] = 34;
// bram[41733] = 20;
// bram[41734] = 10;
// bram[41735] = 3;
// bram[41736] = 0;
// bram[41737] = 0;
// bram[41738] = 5;
// bram[41739] = 12;
// bram[41740] = 24;
// bram[41741] = 38;
// bram[41742] = 55;
// bram[41743] = 74;
// bram[41744] = 95;
// bram[41745] = 117;
// bram[41746] = 138;
// bram[41747] = 160;
// bram[41748] = 181;
// bram[41749] = 200;
// bram[41750] = 216;
// bram[41751] = 230;
// bram[41752] = 241;
// bram[41753] = 249;
// bram[41754] = 253;
// bram[41755] = 253;
// bram[41756] = 250;
// bram[41757] = 242;
// bram[41758] = 232;
// bram[41759] = 218;
// bram[41760] = 201;
// bram[41761] = 182;
// bram[41762] = 162;
// bram[41763] = 140;
// bram[41764] = 119;
// bram[41765] = 97;
// bram[41766] = 76;
// bram[41767] = 57;
// bram[41768] = 40;
// bram[41769] = 25;
// bram[41770] = 13;
// bram[41771] = 5;
// bram[41772] = 1;
// bram[41773] = 0;
// bram[41774] = 3;
// bram[41775] = 9;
// bram[41776] = 19;
// bram[41777] = 33;
// bram[41778] = 49;
// bram[41779] = 67;
// bram[41780] = 87;
// bram[41781] = 109;
// bram[41782] = 130;
// bram[41783] = 152;
// bram[41784] = 173;
// bram[41785] = 193;
// bram[41786] = 210;
// bram[41787] = 226;
// bram[41788] = 238;
// bram[41789] = 247;
// bram[41790] = 252;
// bram[41791] = 253;
// bram[41792] = 251;
// bram[41793] = 245;
// bram[41794] = 236;
// bram[41795] = 223;
// bram[41796] = 207;
// bram[41797] = 189;
// bram[41798] = 170;
// bram[41799] = 148;
// bram[41800] = 126;
// bram[41801] = 105;
// bram[41802] = 83;
// bram[41803] = 64;
// bram[41804] = 46;
// bram[41805] = 30;
// bram[41806] = 17;
// bram[41807] = 8;
// bram[41808] = 2;
// bram[41809] = 0;
// bram[41810] = 1;
// bram[41811] = 6;
// bram[41812] = 15;
// bram[41813] = 27;
// bram[41814] = 43;
// bram[41815] = 60;
// bram[41816] = 80;
// bram[41817] = 101;
// bram[41818] = 123;
// bram[41819] = 144;
// bram[41820] = 166;
// bram[41821] = 186;
// bram[41822] = 204;
// bram[41823] = 220;
// bram[41824] = 234;
// bram[41825] = 244;
// bram[41826] = 250;
// bram[41827] = 253;
// bram[41828] = 252;
// bram[41829] = 248;
// bram[41830] = 240;
// bram[41831] = 228;
// bram[41832] = 213;
// bram[41833] = 196;
// bram[41834] = 177;
// bram[41835] = 156;
// bram[41836] = 134;
// bram[41837] = 113;
// bram[41838] = 91;
// bram[41839] = 71;
// bram[41840] = 52;
// bram[41841] = 35;
// bram[41842] = 21;
// bram[41843] = 11;
// bram[41844] = 3;
// bram[41845] = 0;
// bram[41846] = 0;
// bram[41847] = 4;
// bram[41848] = 12;
// bram[41849] = 23;
// bram[41850] = 37;
// bram[41851] = 53;
// bram[41852] = 72;
// bram[41853] = 93;
// bram[41854] = 115;
// bram[41855] = 136;
// bram[41856] = 158;
// bram[41857] = 179;
// bram[41858] = 198;
// bram[41859] = 215;
// bram[41860] = 229;
// bram[41861] = 241;
// bram[41862] = 248;
// bram[41863] = 253;
// bram[41864] = 253;
// bram[41865] = 250;
// bram[41866] = 243;
// bram[41867] = 233;
// bram[41868] = 219;
// bram[41869] = 203;
// bram[41870] = 184;
// bram[41871] = 164;
// bram[41872] = 142;
// bram[41873] = 121;
// bram[41874] = 99;
// bram[41875] = 78;
// bram[41876] = 58;
// bram[41877] = 41;
// bram[41878] = 26;
// bram[41879] = 14;
// bram[41880] = 6;
// bram[41881] = 1;
// bram[41882] = 0;
// bram[41883] = 2;
// bram[41884] = 8;
// bram[41885] = 18;
// bram[41886] = 31;
// bram[41887] = 47;
// bram[41888] = 65;
// bram[41889] = 85;
// bram[41890] = 107;
// bram[41891] = 128;
// bram[41892] = 150;
// bram[41893] = 171;
// bram[41894] = 191;
// bram[41895] = 209;
// bram[41896] = 224;
// bram[41897] = 237;
// bram[41898] = 246;
// bram[41899] = 252;
// bram[41900] = 254;
// bram[41901] = 252;
// bram[41902] = 246;
// bram[41903] = 237;
// bram[41904] = 224;
// bram[41905] = 209;
// bram[41906] = 191;
// bram[41907] = 171;
// bram[41908] = 150;
// bram[41909] = 128;
// bram[41910] = 107;
// bram[41911] = 85;
// bram[41912] = 65;
// bram[41913] = 47;
// bram[41914] = 31;
// bram[41915] = 18;
// bram[41916] = 8;
// bram[41917] = 2;
// bram[41918] = 0;
// bram[41919] = 1;
// bram[41920] = 6;
// bram[41921] = 14;
// bram[41922] = 26;
// bram[41923] = 41;
// bram[41924] = 58;
// bram[41925] = 78;
// bram[41926] = 99;
// bram[41927] = 121;
// bram[41928] = 142;
// bram[41929] = 164;
// bram[41930] = 184;
// bram[41931] = 203;
// bram[41932] = 219;
// bram[41933] = 233;
// bram[41934] = 243;
// bram[41935] = 250;
// bram[41936] = 253;
// bram[41937] = 253;
// bram[41938] = 248;
// bram[41939] = 241;
// bram[41940] = 229;
// bram[41941] = 215;
// bram[41942] = 198;
// bram[41943] = 179;
// bram[41944] = 158;
// bram[41945] = 136;
// bram[41946] = 115;
// bram[41947] = 93;
// bram[41948] = 72;
// bram[41949] = 53;
// bram[41950] = 37;
// bram[41951] = 23;
// bram[41952] = 12;
// bram[41953] = 4;
// bram[41954] = 0;
// bram[41955] = 0;
// bram[41956] = 3;
// bram[41957] = 11;
// bram[41958] = 21;
// bram[41959] = 35;
// bram[41960] = 52;
// bram[41961] = 71;
// bram[41962] = 91;
// bram[41963] = 113;
// bram[41964] = 134;
// bram[41965] = 156;
// bram[41966] = 177;
// bram[41967] = 196;
// bram[41968] = 213;
// bram[41969] = 228;
// bram[41970] = 240;
// bram[41971] = 248;
// bram[41972] = 252;
// bram[41973] = 253;
// bram[41974] = 250;
// bram[41975] = 244;
// bram[41976] = 234;
// bram[41977] = 220;
// bram[41978] = 204;
// bram[41979] = 186;
// bram[41980] = 166;
// bram[41981] = 144;
// bram[41982] = 123;
// bram[41983] = 101;
// bram[41984] = 80;
// bram[41985] = 60;
// bram[41986] = 43;
// bram[41987] = 27;
// bram[41988] = 15;
// bram[41989] = 6;
// bram[41990] = 1;
// bram[41991] = 0;
// bram[41992] = 2;
// bram[41993] = 8;
// bram[41994] = 17;
// bram[41995] = 30;
// bram[41996] = 46;
// bram[41997] = 64;
// bram[41998] = 83;
// bram[41999] = 105;
// bram[42000] = 127;
// bram[42001] = 148;
// bram[42002] = 170;
// bram[42003] = 189;
// bram[42004] = 207;
// bram[42005] = 223;
// bram[42006] = 236;
// bram[42007] = 245;
// bram[42008] = 251;
// bram[42009] = 253;
// bram[42010] = 252;
// bram[42011] = 247;
// bram[42012] = 238;
// bram[42013] = 226;
// bram[42014] = 210;
// bram[42015] = 193;
// bram[42016] = 173;
// bram[42017] = 152;
// bram[42018] = 130;
// bram[42019] = 109;
// bram[42020] = 87;
// bram[42021] = 67;
// bram[42022] = 49;
// bram[42023] = 33;
// bram[42024] = 19;
// bram[42025] = 9;
// bram[42026] = 3;
// bram[42027] = 0;
// bram[42028] = 1;
// bram[42029] = 5;
// bram[42030] = 13;
// bram[42031] = 25;
// bram[42032] = 40;
// bram[42033] = 57;
// bram[42034] = 76;
// bram[42035] = 97;
// bram[42036] = 119;
// bram[42037] = 140;
// bram[42038] = 162;
// bram[42039] = 182;
// bram[42040] = 201;
// bram[42041] = 218;
// bram[42042] = 232;
// bram[42043] = 242;
// bram[42044] = 250;
// bram[42045] = 253;
// bram[42046] = 253;
// bram[42047] = 249;
// bram[42048] = 241;
// bram[42049] = 230;
// bram[42050] = 216;
// bram[42051] = 200;
// bram[42052] = 181;
// bram[42053] = 160;
// bram[42054] = 138;
// bram[42055] = 117;
// bram[42056] = 95;
// bram[42057] = 74;
// bram[42058] = 55;
// bram[42059] = 38;
// bram[42060] = 24;
// bram[42061] = 12;
// bram[42062] = 5;
// bram[42063] = 0;
// bram[42064] = 0;
// bram[42065] = 3;
// bram[42066] = 10;
// bram[42067] = 20;
// bram[42068] = 34;
// bram[42069] = 50;
// bram[42070] = 69;
// bram[42071] = 89;
// bram[42072] = 111;
// bram[42073] = 132;
// bram[42074] = 154;
// bram[42075] = 175;
// bram[42076] = 195;
// bram[42077] = 212;
// bram[42078] = 227;
// bram[42079] = 239;
// bram[42080] = 247;
// bram[42081] = 252;
// bram[42082] = 253;
// bram[42083] = 251;
// bram[42084] = 245;
// bram[42085] = 235;
// bram[42086] = 222;
// bram[42087] = 206;
// bram[42088] = 188;
// bram[42089] = 168;
// bram[42090] = 146;
// bram[42091] = 125;
// bram[42092] = 103;
// bram[42093] = 82;
// bram[42094] = 62;
// bram[42095] = 44;
// bram[42096] = 29;
// bram[42097] = 16;
// bram[42098] = 7;
// bram[42099] = 1;
// bram[42100] = 0;
// bram[42101] = 1;
// bram[42102] = 7;
// bram[42103] = 16;
// bram[42104] = 29;
// bram[42105] = 44;
// bram[42106] = 62;
// bram[42107] = 82;
// bram[42108] = 103;
// bram[42109] = 125;
// bram[42110] = 146;
// bram[42111] = 168;
// bram[42112] = 188;
// bram[42113] = 206;
// bram[42114] = 222;
// bram[42115] = 235;
// bram[42116] = 245;
// bram[42117] = 251;
// bram[42118] = 253;
// bram[42119] = 252;
// bram[42120] = 247;
// bram[42121] = 239;
// bram[42122] = 227;
// bram[42123] = 212;
// bram[42124] = 195;
// bram[42125] = 175;
// bram[42126] = 154;
// bram[42127] = 132;
// bram[42128] = 111;
// bram[42129] = 89;
// bram[42130] = 69;
// bram[42131] = 50;
// bram[42132] = 34;
// bram[42133] = 20;
// bram[42134] = 10;
// bram[42135] = 3;
// bram[42136] = 0;
// bram[42137] = 0;
// bram[42138] = 5;
// bram[42139] = 12;
// bram[42140] = 24;
// bram[42141] = 38;
// bram[42142] = 55;
// bram[42143] = 74;
// bram[42144] = 95;
// bram[42145] = 117;
// bram[42146] = 138;
// bram[42147] = 160;
// bram[42148] = 181;
// bram[42149] = 200;
// bram[42150] = 216;
// bram[42151] = 230;
// bram[42152] = 241;
// bram[42153] = 249;
// bram[42154] = 253;
// bram[42155] = 253;
// bram[42156] = 250;
// bram[42157] = 242;
// bram[42158] = 232;
// bram[42159] = 218;
// bram[42160] = 201;
// bram[42161] = 182;
// bram[42162] = 162;
// bram[42163] = 140;
// bram[42164] = 119;
// bram[42165] = 97;
// bram[42166] = 76;
// bram[42167] = 57;
// bram[42168] = 40;
// bram[42169] = 25;
// bram[42170] = 13;
// bram[42171] = 5;
// bram[42172] = 1;
// bram[42173] = 0;
// bram[42174] = 3;
// bram[42175] = 9;
// bram[42176] = 19;
// bram[42177] = 33;
// bram[42178] = 49;
// bram[42179] = 67;
// bram[42180] = 87;
// bram[42181] = 109;
// bram[42182] = 130;
// bram[42183] = 152;
// bram[42184] = 173;
// bram[42185] = 193;
// bram[42186] = 210;
// bram[42187] = 226;
// bram[42188] = 238;
// bram[42189] = 247;
// bram[42190] = 252;
// bram[42191] = 253;
// bram[42192] = 251;
// bram[42193] = 245;
// bram[42194] = 236;
// bram[42195] = 223;
// bram[42196] = 207;
// bram[42197] = 189;
// bram[42198] = 170;
// bram[42199] = 148;
// bram[42200] = 126;
// bram[42201] = 105;
// bram[42202] = 83;
// bram[42203] = 64;
// bram[42204] = 46;
// bram[42205] = 30;
// bram[42206] = 17;
// bram[42207] = 8;
// bram[42208] = 2;
// bram[42209] = 0;
// bram[42210] = 1;
// bram[42211] = 6;
// bram[42212] = 15;
// bram[42213] = 27;
// bram[42214] = 43;
// bram[42215] = 60;
// bram[42216] = 80;
// bram[42217] = 101;
// bram[42218] = 123;
// bram[42219] = 144;
// bram[42220] = 166;
// bram[42221] = 186;
// bram[42222] = 204;
// bram[42223] = 220;
// bram[42224] = 234;
// bram[42225] = 244;
// bram[42226] = 250;
// bram[42227] = 253;
// bram[42228] = 252;
// bram[42229] = 248;
// bram[42230] = 240;
// bram[42231] = 228;
// bram[42232] = 213;
// bram[42233] = 196;
// bram[42234] = 177;
// bram[42235] = 156;
// bram[42236] = 134;
// bram[42237] = 113;
// bram[42238] = 91;
// bram[42239] = 71;
// bram[42240] = 52;
// bram[42241] = 35;
// bram[42242] = 21;
// bram[42243] = 11;
// bram[42244] = 3;
// bram[42245] = 0;
// bram[42246] = 0;
// bram[42247] = 4;
// bram[42248] = 12;
// bram[42249] = 23;
// bram[42250] = 37;
// bram[42251] = 53;
// bram[42252] = 72;
// bram[42253] = 93;
// bram[42254] = 115;
// bram[42255] = 136;
// bram[42256] = 158;
// bram[42257] = 179;
// bram[42258] = 198;
// bram[42259] = 215;
// bram[42260] = 229;
// bram[42261] = 241;
// bram[42262] = 248;
// bram[42263] = 253;
// bram[42264] = 253;
// bram[42265] = 250;
// bram[42266] = 243;
// bram[42267] = 233;
// bram[42268] = 219;
// bram[42269] = 203;
// bram[42270] = 184;
// bram[42271] = 164;
// bram[42272] = 142;
// bram[42273] = 121;
// bram[42274] = 99;
// bram[42275] = 78;
// bram[42276] = 58;
// bram[42277] = 41;
// bram[42278] = 26;
// bram[42279] = 14;
// bram[42280] = 6;
// bram[42281] = 1;
// bram[42282] = 0;
// bram[42283] = 2;
// bram[42284] = 8;
// bram[42285] = 18;
// bram[42286] = 31;
// bram[42287] = 47;
// bram[42288] = 65;
// bram[42289] = 85;
// bram[42290] = 107;
// bram[42291] = 128;
// bram[42292] = 150;
// bram[42293] = 171;
// bram[42294] = 191;
// bram[42295] = 209;
// bram[42296] = 224;
// bram[42297] = 237;
// bram[42298] = 246;
// bram[42299] = 252;
// bram[42300] = 254;
// bram[42301] = 252;
// bram[42302] = 246;
// bram[42303] = 237;
// bram[42304] = 224;
// bram[42305] = 209;
// bram[42306] = 191;
// bram[42307] = 171;
// bram[42308] = 150;
// bram[42309] = 128;
// bram[42310] = 107;
// bram[42311] = 85;
// bram[42312] = 65;
// bram[42313] = 47;
// bram[42314] = 31;
// bram[42315] = 18;
// bram[42316] = 8;
// bram[42317] = 2;
// bram[42318] = 0;
// bram[42319] = 1;
// bram[42320] = 6;
// bram[42321] = 14;
// bram[42322] = 26;
// bram[42323] = 41;
// bram[42324] = 58;
// bram[42325] = 78;
// bram[42326] = 99;
// bram[42327] = 121;
// bram[42328] = 142;
// bram[42329] = 164;
// bram[42330] = 184;
// bram[42331] = 203;
// bram[42332] = 219;
// bram[42333] = 233;
// bram[42334] = 243;
// bram[42335] = 250;
// bram[42336] = 253;
// bram[42337] = 253;
// bram[42338] = 248;
// bram[42339] = 241;
// bram[42340] = 229;
// bram[42341] = 215;
// bram[42342] = 198;
// bram[42343] = 179;
// bram[42344] = 158;
// bram[42345] = 136;
// bram[42346] = 115;
// bram[42347] = 93;
// bram[42348] = 72;
// bram[42349] = 53;
// bram[42350] = 37;
// bram[42351] = 23;
// bram[42352] = 12;
// bram[42353] = 4;
// bram[42354] = 0;
// bram[42355] = 0;
// bram[42356] = 3;
// bram[42357] = 11;
// bram[42358] = 21;
// bram[42359] = 35;
// bram[42360] = 52;
// bram[42361] = 71;
// bram[42362] = 91;
// bram[42363] = 113;
// bram[42364] = 134;
// bram[42365] = 156;
// bram[42366] = 177;
// bram[42367] = 196;
// bram[42368] = 213;
// bram[42369] = 228;
// bram[42370] = 240;
// bram[42371] = 248;
// bram[42372] = 252;
// bram[42373] = 253;
// bram[42374] = 250;
// bram[42375] = 244;
// bram[42376] = 234;
// bram[42377] = 220;
// bram[42378] = 204;
// bram[42379] = 186;
// bram[42380] = 166;
// bram[42381] = 144;
// bram[42382] = 123;
// bram[42383] = 101;
// bram[42384] = 80;
// bram[42385] = 60;
// bram[42386] = 43;
// bram[42387] = 27;
// bram[42388] = 15;
// bram[42389] = 6;
// bram[42390] = 1;
// bram[42391] = 0;
// bram[42392] = 2;
// bram[42393] = 8;
// bram[42394] = 17;
// bram[42395] = 30;
// bram[42396] = 46;
// bram[42397] = 64;
// bram[42398] = 83;
// bram[42399] = 105;
// bram[42400] = 126;
// bram[42401] = 148;
// bram[42402] = 170;
// bram[42403] = 189;
// bram[42404] = 207;
// bram[42405] = 223;
// bram[42406] = 236;
// bram[42407] = 245;
// bram[42408] = 251;
// bram[42409] = 253;
// bram[42410] = 252;
// bram[42411] = 247;
// bram[42412] = 238;
// bram[42413] = 226;
// bram[42414] = 210;
// bram[42415] = 193;
// bram[42416] = 173;
// bram[42417] = 152;
// bram[42418] = 130;
// bram[42419] = 109;
// bram[42420] = 87;
// bram[42421] = 67;
// bram[42422] = 49;
// bram[42423] = 33;
// bram[42424] = 19;
// bram[42425] = 9;
// bram[42426] = 3;
// bram[42427] = 0;
// bram[42428] = 1;
// bram[42429] = 5;
// bram[42430] = 13;
// bram[42431] = 25;
// bram[42432] = 40;
// bram[42433] = 57;
// bram[42434] = 76;
// bram[42435] = 97;
// bram[42436] = 119;
// bram[42437] = 140;
// bram[42438] = 162;
// bram[42439] = 182;
// bram[42440] = 201;
// bram[42441] = 218;
// bram[42442] = 232;
// bram[42443] = 242;
// bram[42444] = 250;
// bram[42445] = 253;
// bram[42446] = 253;
// bram[42447] = 249;
// bram[42448] = 241;
// bram[42449] = 230;
// bram[42450] = 216;
// bram[42451] = 200;
// bram[42452] = 181;
// bram[42453] = 160;
// bram[42454] = 138;
// bram[42455] = 117;
// bram[42456] = 95;
// bram[42457] = 74;
// bram[42458] = 55;
// bram[42459] = 38;
// bram[42460] = 24;
// bram[42461] = 12;
// bram[42462] = 5;
// bram[42463] = 0;
// bram[42464] = 0;
// bram[42465] = 3;
// bram[42466] = 10;
// bram[42467] = 20;
// bram[42468] = 34;
// bram[42469] = 50;
// bram[42470] = 69;
// bram[42471] = 89;
// bram[42472] = 111;
// bram[42473] = 132;
// bram[42474] = 154;
// bram[42475] = 175;
// bram[42476] = 195;
// bram[42477] = 212;
// bram[42478] = 227;
// bram[42479] = 239;
// bram[42480] = 247;
// bram[42481] = 252;
// bram[42482] = 253;
// bram[42483] = 251;
// bram[42484] = 245;
// bram[42485] = 235;
// bram[42486] = 222;
// bram[42487] = 206;
// bram[42488] = 188;
// bram[42489] = 168;
// bram[42490] = 146;
// bram[42491] = 125;
// bram[42492] = 103;
// bram[42493] = 82;
// bram[42494] = 62;
// bram[42495] = 44;
// bram[42496] = 29;
// bram[42497] = 16;
// bram[42498] = 7;
// bram[42499] = 1;
// bram[42500] = 0;
// bram[42501] = 1;
// bram[42502] = 7;
// bram[42503] = 16;
// bram[42504] = 29;
// bram[42505] = 44;
// bram[42506] = 62;
// bram[42507] = 82;
// bram[42508] = 103;
// bram[42509] = 125;
// bram[42510] = 146;
// bram[42511] = 168;
// bram[42512] = 188;
// bram[42513] = 206;
// bram[42514] = 222;
// bram[42515] = 235;
// bram[42516] = 245;
// bram[42517] = 251;
// bram[42518] = 253;
// bram[42519] = 252;
// bram[42520] = 247;
// bram[42521] = 239;
// bram[42522] = 227;
// bram[42523] = 212;
// bram[42524] = 195;
// bram[42525] = 175;
// bram[42526] = 154;
// bram[42527] = 132;
// bram[42528] = 111;
// bram[42529] = 89;
// bram[42530] = 69;
// bram[42531] = 50;
// bram[42532] = 34;
// bram[42533] = 20;
// bram[42534] = 10;
// bram[42535] = 3;
// bram[42536] = 0;
// bram[42537] = 0;
// bram[42538] = 5;
// bram[42539] = 12;
// bram[42540] = 24;
// bram[42541] = 38;
// bram[42542] = 55;
// bram[42543] = 74;
// bram[42544] = 95;
// bram[42545] = 117;
// bram[42546] = 138;
// bram[42547] = 160;
// bram[42548] = 181;
// bram[42549] = 200;
// bram[42550] = 216;
// bram[42551] = 230;
// bram[42552] = 241;
// bram[42553] = 249;
// bram[42554] = 253;
// bram[42555] = 253;
// bram[42556] = 250;
// bram[42557] = 242;
// bram[42558] = 232;
// bram[42559] = 218;
// bram[42560] = 201;
// bram[42561] = 182;
// bram[42562] = 162;
// bram[42563] = 140;
// bram[42564] = 119;
// bram[42565] = 97;
// bram[42566] = 76;
// bram[42567] = 57;
// bram[42568] = 40;
// bram[42569] = 25;
// bram[42570] = 13;
// bram[42571] = 5;
// bram[42572] = 1;
// bram[42573] = 0;
// bram[42574] = 3;
// bram[42575] = 9;
// bram[42576] = 19;
// bram[42577] = 33;
// bram[42578] = 49;
// bram[42579] = 67;
// bram[42580] = 87;
// bram[42581] = 109;
// bram[42582] = 130;
// bram[42583] = 152;
// bram[42584] = 173;
// bram[42585] = 193;
// bram[42586] = 210;
// bram[42587] = 226;
// bram[42588] = 238;
// bram[42589] = 247;
// bram[42590] = 252;
// bram[42591] = 253;
// bram[42592] = 251;
// bram[42593] = 245;
// bram[42594] = 236;
// bram[42595] = 223;
// bram[42596] = 207;
// bram[42597] = 189;
// bram[42598] = 170;
// bram[42599] = 148;
// bram[42600] = 126;
// bram[42601] = 105;
// bram[42602] = 83;
// bram[42603] = 64;
// bram[42604] = 46;
// bram[42605] = 30;
// bram[42606] = 17;
// bram[42607] = 8;
// bram[42608] = 2;
// bram[42609] = 0;
// bram[42610] = 1;
// bram[42611] = 6;
// bram[42612] = 15;
// bram[42613] = 27;
// bram[42614] = 43;
// bram[42615] = 60;
// bram[42616] = 80;
// bram[42617] = 101;
// bram[42618] = 123;
// bram[42619] = 144;
// bram[42620] = 166;
// bram[42621] = 186;
// bram[42622] = 204;
// bram[42623] = 220;
// bram[42624] = 234;
// bram[42625] = 244;
// bram[42626] = 250;
// bram[42627] = 253;
// bram[42628] = 252;
// bram[42629] = 248;
// bram[42630] = 240;
// bram[42631] = 228;
// bram[42632] = 213;
// bram[42633] = 196;
// bram[42634] = 177;
// bram[42635] = 156;
// bram[42636] = 134;
// bram[42637] = 113;
// bram[42638] = 91;
// bram[42639] = 71;
// bram[42640] = 52;
// bram[42641] = 35;
// bram[42642] = 21;
// bram[42643] = 11;
// bram[42644] = 3;
// bram[42645] = 0;
// bram[42646] = 0;
// bram[42647] = 4;
// bram[42648] = 12;
// bram[42649] = 23;
// bram[42650] = 37;
// bram[42651] = 53;
// bram[42652] = 72;
// bram[42653] = 93;
// bram[42654] = 115;
// bram[42655] = 136;
// bram[42656] = 158;
// bram[42657] = 179;
// bram[42658] = 198;
// bram[42659] = 215;
// bram[42660] = 229;
// bram[42661] = 241;
// bram[42662] = 248;
// bram[42663] = 253;
// bram[42664] = 253;
// bram[42665] = 250;
// bram[42666] = 243;
// bram[42667] = 233;
// bram[42668] = 219;
// bram[42669] = 203;
// bram[42670] = 184;
// bram[42671] = 164;
// bram[42672] = 142;
// bram[42673] = 121;
// bram[42674] = 99;
// bram[42675] = 78;
// bram[42676] = 58;
// bram[42677] = 41;
// bram[42678] = 26;
// bram[42679] = 14;
// bram[42680] = 6;
// bram[42681] = 1;
// bram[42682] = 0;
// bram[42683] = 2;
// bram[42684] = 8;
// bram[42685] = 18;
// bram[42686] = 31;
// bram[42687] = 47;
// bram[42688] = 65;
// bram[42689] = 85;
// bram[42690] = 107;
// bram[42691] = 128;
// bram[42692] = 150;
// bram[42693] = 171;
// bram[42694] = 191;
// bram[42695] = 209;
// bram[42696] = 224;
// bram[42697] = 237;
// bram[42698] = 246;
// bram[42699] = 252;
// bram[42700] = 254;
// bram[42701] = 252;
// bram[42702] = 246;
// bram[42703] = 237;
// bram[42704] = 224;
// bram[42705] = 209;
// bram[42706] = 191;
// bram[42707] = 171;
// bram[42708] = 150;
// bram[42709] = 128;
// bram[42710] = 107;
// bram[42711] = 85;
// bram[42712] = 65;
// bram[42713] = 47;
// bram[42714] = 31;
// bram[42715] = 18;
// bram[42716] = 8;
// bram[42717] = 2;
// bram[42718] = 0;
// bram[42719] = 1;
// bram[42720] = 6;
// bram[42721] = 14;
// bram[42722] = 26;
// bram[42723] = 41;
// bram[42724] = 58;
// bram[42725] = 78;
// bram[42726] = 99;
// bram[42727] = 121;
// bram[42728] = 142;
// bram[42729] = 164;
// bram[42730] = 184;
// bram[42731] = 203;
// bram[42732] = 219;
// bram[42733] = 233;
// bram[42734] = 243;
// bram[42735] = 250;
// bram[42736] = 253;
// bram[42737] = 253;
// bram[42738] = 248;
// bram[42739] = 241;
// bram[42740] = 229;
// bram[42741] = 215;
// bram[42742] = 198;
// bram[42743] = 179;
// bram[42744] = 158;
// bram[42745] = 136;
// bram[42746] = 115;
// bram[42747] = 93;
// bram[42748] = 72;
// bram[42749] = 53;
// bram[42750] = 37;
// bram[42751] = 23;
// bram[42752] = 12;
// bram[42753] = 4;
// bram[42754] = 0;
// bram[42755] = 0;
// bram[42756] = 3;
// bram[42757] = 11;
// bram[42758] = 21;
// bram[42759] = 35;
// bram[42760] = 52;
// bram[42761] = 71;
// bram[42762] = 91;
// bram[42763] = 113;
// bram[42764] = 134;
// bram[42765] = 156;
// bram[42766] = 177;
// bram[42767] = 196;
// bram[42768] = 213;
// bram[42769] = 228;
// bram[42770] = 240;
// bram[42771] = 248;
// bram[42772] = 252;
// bram[42773] = 253;
// bram[42774] = 250;
// bram[42775] = 244;
// bram[42776] = 234;
// bram[42777] = 220;
// bram[42778] = 204;
// bram[42779] = 186;
// bram[42780] = 166;
// bram[42781] = 144;
// bram[42782] = 123;
// bram[42783] = 101;
// bram[42784] = 80;
// bram[42785] = 60;
// bram[42786] = 43;
// bram[42787] = 27;
// bram[42788] = 15;
// bram[42789] = 6;
// bram[42790] = 1;
// bram[42791] = 0;
// bram[42792] = 2;
// bram[42793] = 8;
// bram[42794] = 17;
// bram[42795] = 30;
// bram[42796] = 46;
// bram[42797] = 64;
// bram[42798] = 83;
// bram[42799] = 105;
// bram[42800] = 127;
// bram[42801] = 148;
// bram[42802] = 170;
// bram[42803] = 189;
// bram[42804] = 207;
// bram[42805] = 223;
// bram[42806] = 236;
// bram[42807] = 245;
// bram[42808] = 251;
// bram[42809] = 253;
// bram[42810] = 252;
// bram[42811] = 247;
// bram[42812] = 238;
// bram[42813] = 226;
// bram[42814] = 210;
// bram[42815] = 193;
// bram[42816] = 173;
// bram[42817] = 152;
// bram[42818] = 130;
// bram[42819] = 109;
// bram[42820] = 87;
// bram[42821] = 67;
// bram[42822] = 49;
// bram[42823] = 33;
// bram[42824] = 19;
// bram[42825] = 9;
// bram[42826] = 3;
// bram[42827] = 0;
// bram[42828] = 1;
// bram[42829] = 5;
// bram[42830] = 13;
// bram[42831] = 25;
// bram[42832] = 40;
// bram[42833] = 57;
// bram[42834] = 76;
// bram[42835] = 97;
// bram[42836] = 119;
// bram[42837] = 140;
// bram[42838] = 162;
// bram[42839] = 182;
// bram[42840] = 201;
// bram[42841] = 218;
// bram[42842] = 232;
// bram[42843] = 242;
// bram[42844] = 250;
// bram[42845] = 253;
// bram[42846] = 253;
// bram[42847] = 249;
// bram[42848] = 241;
// bram[42849] = 230;
// bram[42850] = 216;
// bram[42851] = 200;
// bram[42852] = 181;
// bram[42853] = 160;
// bram[42854] = 138;
// bram[42855] = 117;
// bram[42856] = 95;
// bram[42857] = 74;
// bram[42858] = 55;
// bram[42859] = 38;
// bram[42860] = 24;
// bram[42861] = 12;
// bram[42862] = 5;
// bram[42863] = 0;
// bram[42864] = 0;
// bram[42865] = 3;
// bram[42866] = 10;
// bram[42867] = 20;
// bram[42868] = 34;
// bram[42869] = 50;
// bram[42870] = 69;
// bram[42871] = 89;
// bram[42872] = 111;
// bram[42873] = 132;
// bram[42874] = 154;
// bram[42875] = 175;
// bram[42876] = 195;
// bram[42877] = 212;
// bram[42878] = 227;
// bram[42879] = 239;
// bram[42880] = 247;
// bram[42881] = 252;
// bram[42882] = 253;
// bram[42883] = 251;
// bram[42884] = 245;
// bram[42885] = 235;
// bram[42886] = 222;
// bram[42887] = 206;
// bram[42888] = 188;
// bram[42889] = 168;
// bram[42890] = 146;
// bram[42891] = 125;
// bram[42892] = 103;
// bram[42893] = 82;
// bram[42894] = 62;
// bram[42895] = 44;
// bram[42896] = 29;
// bram[42897] = 16;
// bram[42898] = 7;
// bram[42899] = 1;
// bram[42900] = 0;
// bram[42901] = 1;
// bram[42902] = 7;
// bram[42903] = 16;
// bram[42904] = 29;
// bram[42905] = 44;
// bram[42906] = 62;
// bram[42907] = 82;
// bram[42908] = 103;
// bram[42909] = 125;
// bram[42910] = 146;
// bram[42911] = 168;
// bram[42912] = 188;
// bram[42913] = 206;
// bram[42914] = 222;
// bram[42915] = 235;
// bram[42916] = 245;
// bram[42917] = 251;
// bram[42918] = 253;
// bram[42919] = 252;
// bram[42920] = 247;
// bram[42921] = 239;
// bram[42922] = 227;
// bram[42923] = 212;
// bram[42924] = 195;
// bram[42925] = 175;
// bram[42926] = 154;
// bram[42927] = 132;
// bram[42928] = 111;
// bram[42929] = 89;
// bram[42930] = 69;
// bram[42931] = 50;
// bram[42932] = 34;
// bram[42933] = 20;
// bram[42934] = 10;
// bram[42935] = 3;
// bram[42936] = 0;
// bram[42937] = 0;
// bram[42938] = 5;
// bram[42939] = 12;
// bram[42940] = 24;
// bram[42941] = 38;
// bram[42942] = 55;
// bram[42943] = 74;
// bram[42944] = 95;
// bram[42945] = 117;
// bram[42946] = 138;
// bram[42947] = 160;
// bram[42948] = 181;
// bram[42949] = 200;
// bram[42950] = 216;
// bram[42951] = 230;
// bram[42952] = 241;
// bram[42953] = 249;
// bram[42954] = 253;
// bram[42955] = 253;
// bram[42956] = 250;
// bram[42957] = 242;
// bram[42958] = 232;
// bram[42959] = 218;
// bram[42960] = 201;
// bram[42961] = 182;
// bram[42962] = 162;
// bram[42963] = 140;
// bram[42964] = 119;
// bram[42965] = 97;
// bram[42966] = 76;
// bram[42967] = 57;
// bram[42968] = 40;
// bram[42969] = 25;
// bram[42970] = 13;
// bram[42971] = 5;
// bram[42972] = 1;
// bram[42973] = 0;
// bram[42974] = 3;
// bram[42975] = 9;
// bram[42976] = 19;
// bram[42977] = 33;
// bram[42978] = 49;
// bram[42979] = 67;
// bram[42980] = 87;
// bram[42981] = 109;
// bram[42982] = 130;
// bram[42983] = 152;
// bram[42984] = 173;
// bram[42985] = 193;
// bram[42986] = 210;
// bram[42987] = 226;
// bram[42988] = 238;
// bram[42989] = 247;
// bram[42990] = 252;
// bram[42991] = 253;
// bram[42992] = 251;
// bram[42993] = 245;
// bram[42994] = 236;
// bram[42995] = 223;
// bram[42996] = 207;
// bram[42997] = 189;
// bram[42998] = 170;
// bram[42999] = 148;
// bram[43000] = 126;
// bram[43001] = 105;
// bram[43002] = 83;
// bram[43003] = 64;
// bram[43004] = 46;
// bram[43005] = 30;
// bram[43006] = 17;
// bram[43007] = 8;
// bram[43008] = 2;
// bram[43009] = 0;
// bram[43010] = 1;
// bram[43011] = 6;
// bram[43012] = 15;
// bram[43013] = 27;
// bram[43014] = 43;
// bram[43015] = 60;
// bram[43016] = 80;
// bram[43017] = 101;
// bram[43018] = 123;
// bram[43019] = 144;
// bram[43020] = 166;
// bram[43021] = 186;
// bram[43022] = 204;
// bram[43023] = 220;
// bram[43024] = 234;
// bram[43025] = 244;
// bram[43026] = 250;
// bram[43027] = 253;
// bram[43028] = 252;
// bram[43029] = 248;
// bram[43030] = 240;
// bram[43031] = 228;
// bram[43032] = 213;
// bram[43033] = 196;
// bram[43034] = 177;
// bram[43035] = 156;
// bram[43036] = 134;
// bram[43037] = 113;
// bram[43038] = 91;
// bram[43039] = 71;
// bram[43040] = 52;
// bram[43041] = 35;
// bram[43042] = 21;
// bram[43043] = 11;
// bram[43044] = 3;
// bram[43045] = 0;
// bram[43046] = 0;
// bram[43047] = 4;
// bram[43048] = 12;
// bram[43049] = 23;
// bram[43050] = 37;
// bram[43051] = 53;
// bram[43052] = 72;
// bram[43053] = 93;
// bram[43054] = 115;
// bram[43055] = 136;
// bram[43056] = 158;
// bram[43057] = 179;
// bram[43058] = 198;
// bram[43059] = 215;
// bram[43060] = 229;
// bram[43061] = 241;
// bram[43062] = 248;
// bram[43063] = 253;
// bram[43064] = 253;
// bram[43065] = 250;
// bram[43066] = 243;
// bram[43067] = 233;
// bram[43068] = 219;
// bram[43069] = 203;
// bram[43070] = 184;
// bram[43071] = 164;
// bram[43072] = 142;
// bram[43073] = 121;
// bram[43074] = 99;
// bram[43075] = 78;
// bram[43076] = 58;
// bram[43077] = 41;
// bram[43078] = 26;
// bram[43079] = 14;
// bram[43080] = 6;
// bram[43081] = 1;
// bram[43082] = 0;
// bram[43083] = 2;
// bram[43084] = 8;
// bram[43085] = 18;
// bram[43086] = 31;
// bram[43087] = 47;
// bram[43088] = 65;
// bram[43089] = 85;
// bram[43090] = 107;
// bram[43091] = 128;
// bram[43092] = 150;
// bram[43093] = 171;
// bram[43094] = 191;
// bram[43095] = 209;
// bram[43096] = 224;
// bram[43097] = 237;
// bram[43098] = 246;
// bram[43099] = 252;
// bram[43100] = 254;
// bram[43101] = 252;
// bram[43102] = 246;
// bram[43103] = 237;
// bram[43104] = 224;
// bram[43105] = 209;
// bram[43106] = 191;
// bram[43107] = 171;
// bram[43108] = 150;
// bram[43109] = 128;
// bram[43110] = 107;
// bram[43111] = 85;
// bram[43112] = 65;
// bram[43113] = 47;
// bram[43114] = 31;
// bram[43115] = 18;
// bram[43116] = 8;
// bram[43117] = 2;
// bram[43118] = 0;
// bram[43119] = 1;
// bram[43120] = 6;
// bram[43121] = 14;
// bram[43122] = 26;
// bram[43123] = 41;
// bram[43124] = 58;
// bram[43125] = 78;
// bram[43126] = 99;
// bram[43127] = 121;
// bram[43128] = 142;
// bram[43129] = 164;
// bram[43130] = 184;
// bram[43131] = 203;
// bram[43132] = 219;
// bram[43133] = 233;
// bram[43134] = 243;
// bram[43135] = 250;
// bram[43136] = 253;
// bram[43137] = 253;
// bram[43138] = 248;
// bram[43139] = 241;
// bram[43140] = 229;
// bram[43141] = 215;
// bram[43142] = 198;
// bram[43143] = 179;
// bram[43144] = 158;
// bram[43145] = 136;
// bram[43146] = 115;
// bram[43147] = 93;
// bram[43148] = 72;
// bram[43149] = 53;
// bram[43150] = 37;
// bram[43151] = 23;
// bram[43152] = 12;
// bram[43153] = 4;
// bram[43154] = 0;
// bram[43155] = 0;
// bram[43156] = 3;
// bram[43157] = 11;
// bram[43158] = 21;
// bram[43159] = 35;
// bram[43160] = 52;
// bram[43161] = 71;
// bram[43162] = 91;
// bram[43163] = 113;
// bram[43164] = 134;
// bram[43165] = 156;
// bram[43166] = 177;
// bram[43167] = 196;
// bram[43168] = 213;
// bram[43169] = 228;
// bram[43170] = 240;
// bram[43171] = 248;
// bram[43172] = 252;
// bram[43173] = 253;
// bram[43174] = 250;
// bram[43175] = 244;
// bram[43176] = 234;
// bram[43177] = 220;
// bram[43178] = 204;
// bram[43179] = 186;
// bram[43180] = 166;
// bram[43181] = 144;
// bram[43182] = 123;
// bram[43183] = 101;
// bram[43184] = 80;
// bram[43185] = 60;
// bram[43186] = 43;
// bram[43187] = 27;
// bram[43188] = 15;
// bram[43189] = 6;
// bram[43190] = 1;
// bram[43191] = 0;
// bram[43192] = 2;
// bram[43193] = 8;
// bram[43194] = 17;
// bram[43195] = 30;
// bram[43196] = 46;
// bram[43197] = 64;
// bram[43198] = 83;
// bram[43199] = 105;
// bram[43200] = 127;
// bram[43201] = 148;
// bram[43202] = 170;
// bram[43203] = 189;
// bram[43204] = 207;
// bram[43205] = 223;
// bram[43206] = 236;
// bram[43207] = 245;
// bram[43208] = 251;
// bram[43209] = 253;
// bram[43210] = 252;
// bram[43211] = 247;
// bram[43212] = 238;
// bram[43213] = 226;
// bram[43214] = 210;
// bram[43215] = 193;
// bram[43216] = 173;
// bram[43217] = 152;
// bram[43218] = 130;
// bram[43219] = 109;
// bram[43220] = 87;
// bram[43221] = 67;
// bram[43222] = 49;
// bram[43223] = 33;
// bram[43224] = 19;
// bram[43225] = 9;
// bram[43226] = 3;
// bram[43227] = 0;
// bram[43228] = 1;
// bram[43229] = 5;
// bram[43230] = 13;
// bram[43231] = 25;
// bram[43232] = 40;
// bram[43233] = 57;
// bram[43234] = 76;
// bram[43235] = 97;
// bram[43236] = 119;
// bram[43237] = 140;
// bram[43238] = 162;
// bram[43239] = 182;
// bram[43240] = 201;
// bram[43241] = 218;
// bram[43242] = 232;
// bram[43243] = 242;
// bram[43244] = 250;
// bram[43245] = 253;
// bram[43246] = 253;
// bram[43247] = 249;
// bram[43248] = 241;
// bram[43249] = 230;
// bram[43250] = 216;
// bram[43251] = 200;
// bram[43252] = 181;
// bram[43253] = 160;
// bram[43254] = 138;
// bram[43255] = 117;
// bram[43256] = 95;
// bram[43257] = 74;
// bram[43258] = 55;
// bram[43259] = 38;
// bram[43260] = 24;
// bram[43261] = 12;
// bram[43262] = 5;
// bram[43263] = 0;
// bram[43264] = 0;
// bram[43265] = 3;
// bram[43266] = 10;
// bram[43267] = 20;
// bram[43268] = 34;
// bram[43269] = 50;
// bram[43270] = 69;
// bram[43271] = 89;
// bram[43272] = 111;
// bram[43273] = 132;
// bram[43274] = 154;
// bram[43275] = 175;
// bram[43276] = 195;
// bram[43277] = 212;
// bram[43278] = 227;
// bram[43279] = 239;
// bram[43280] = 247;
// bram[43281] = 252;
// bram[43282] = 253;
// bram[43283] = 251;
// bram[43284] = 245;
// bram[43285] = 235;
// bram[43286] = 222;
// bram[43287] = 206;
// bram[43288] = 188;
// bram[43289] = 168;
// bram[43290] = 146;
// bram[43291] = 125;
// bram[43292] = 103;
// bram[43293] = 82;
// bram[43294] = 62;
// bram[43295] = 44;
// bram[43296] = 29;
// bram[43297] = 16;
// bram[43298] = 7;
// bram[43299] = 1;
// bram[43300] = 0;
// bram[43301] = 1;
// bram[43302] = 7;
// bram[43303] = 16;
// bram[43304] = 29;
// bram[43305] = 44;
// bram[43306] = 62;
// bram[43307] = 82;
// bram[43308] = 103;
// bram[43309] = 125;
// bram[43310] = 146;
// bram[43311] = 168;
// bram[43312] = 188;
// bram[43313] = 206;
// bram[43314] = 222;
// bram[43315] = 235;
// bram[43316] = 245;
// bram[43317] = 251;
// bram[43318] = 253;
// bram[43319] = 252;
// bram[43320] = 247;
// bram[43321] = 239;
// bram[43322] = 227;
// bram[43323] = 212;
// bram[43324] = 195;
// bram[43325] = 175;
// bram[43326] = 154;
// bram[43327] = 132;
// bram[43328] = 111;
// bram[43329] = 89;
// bram[43330] = 69;
// bram[43331] = 50;
// bram[43332] = 34;
// bram[43333] = 20;
// bram[43334] = 10;
// bram[43335] = 3;
// bram[43336] = 0;
// bram[43337] = 0;
// bram[43338] = 5;
// bram[43339] = 12;
// bram[43340] = 24;
// bram[43341] = 38;
// bram[43342] = 55;
// bram[43343] = 74;
// bram[43344] = 95;
// bram[43345] = 117;
// bram[43346] = 138;
// bram[43347] = 160;
// bram[43348] = 181;
// bram[43349] = 200;
// bram[43350] = 216;
// bram[43351] = 230;
// bram[43352] = 241;
// bram[43353] = 249;
// bram[43354] = 253;
// bram[43355] = 253;
// bram[43356] = 250;
// bram[43357] = 242;
// bram[43358] = 232;
// bram[43359] = 218;
// bram[43360] = 201;
// bram[43361] = 182;
// bram[43362] = 162;
// bram[43363] = 140;
// bram[43364] = 119;
// bram[43365] = 97;
// bram[43366] = 76;
// bram[43367] = 57;
// bram[43368] = 40;
// bram[43369] = 25;
// bram[43370] = 13;
// bram[43371] = 5;
// bram[43372] = 1;
// bram[43373] = 0;
// bram[43374] = 3;
// bram[43375] = 9;
// bram[43376] = 19;
// bram[43377] = 33;
// bram[43378] = 49;
// bram[43379] = 67;
// bram[43380] = 87;
// bram[43381] = 109;
// bram[43382] = 130;
// bram[43383] = 152;
// bram[43384] = 173;
// bram[43385] = 193;
// bram[43386] = 210;
// bram[43387] = 226;
// bram[43388] = 238;
// bram[43389] = 247;
// bram[43390] = 252;
// bram[43391] = 253;
// bram[43392] = 251;
// bram[43393] = 245;
// bram[43394] = 236;
// bram[43395] = 223;
// bram[43396] = 207;
// bram[43397] = 189;
// bram[43398] = 170;
// bram[43399] = 148;
// bram[43400] = 126;
// bram[43401] = 105;
// bram[43402] = 83;
// bram[43403] = 64;
// bram[43404] = 46;
// bram[43405] = 30;
// bram[43406] = 17;
// bram[43407] = 8;
// bram[43408] = 2;
// bram[43409] = 0;
// bram[43410] = 1;
// bram[43411] = 6;
// bram[43412] = 15;
// bram[43413] = 27;
// bram[43414] = 43;
// bram[43415] = 60;
// bram[43416] = 80;
// bram[43417] = 101;
// bram[43418] = 123;
// bram[43419] = 144;
// bram[43420] = 166;
// bram[43421] = 186;
// bram[43422] = 204;
// bram[43423] = 220;
// bram[43424] = 234;
// bram[43425] = 244;
// bram[43426] = 250;
// bram[43427] = 253;
// bram[43428] = 252;
// bram[43429] = 248;
// bram[43430] = 240;
// bram[43431] = 228;
// bram[43432] = 213;
// bram[43433] = 196;
// bram[43434] = 177;
// bram[43435] = 156;
// bram[43436] = 134;
// bram[43437] = 113;
// bram[43438] = 91;
// bram[43439] = 71;
// bram[43440] = 52;
// bram[43441] = 35;
// bram[43442] = 21;
// bram[43443] = 11;
// bram[43444] = 3;
// bram[43445] = 0;
// bram[43446] = 0;
// bram[43447] = 4;
// bram[43448] = 12;
// bram[43449] = 23;
// bram[43450] = 37;
// bram[43451] = 53;
// bram[43452] = 72;
// bram[43453] = 93;
// bram[43454] = 115;
// bram[43455] = 136;
// bram[43456] = 158;
// bram[43457] = 179;
// bram[43458] = 198;
// bram[43459] = 215;
// bram[43460] = 229;
// bram[43461] = 241;
// bram[43462] = 248;
// bram[43463] = 253;
// bram[43464] = 253;
// bram[43465] = 250;
// bram[43466] = 243;
// bram[43467] = 233;
// bram[43468] = 219;
// bram[43469] = 203;
// bram[43470] = 184;
// bram[43471] = 164;
// bram[43472] = 142;
// bram[43473] = 121;
// bram[43474] = 99;
// bram[43475] = 78;
// bram[43476] = 58;
// bram[43477] = 41;
// bram[43478] = 26;
// bram[43479] = 14;
// bram[43480] = 6;
// bram[43481] = 1;
// bram[43482] = 0;
// bram[43483] = 2;
// bram[43484] = 8;
// bram[43485] = 18;
// bram[43486] = 31;
// bram[43487] = 47;
// bram[43488] = 65;
// bram[43489] = 85;
// bram[43490] = 107;
// bram[43491] = 128;
// bram[43492] = 150;
// bram[43493] = 171;
// bram[43494] = 191;
// bram[43495] = 209;
// bram[43496] = 224;
// bram[43497] = 237;
// bram[43498] = 246;
// bram[43499] = 252;
// bram[43500] = 254;
// bram[43501] = 252;
// bram[43502] = 246;
// bram[43503] = 237;
// bram[43504] = 224;
// bram[43505] = 209;
// bram[43506] = 191;
// bram[43507] = 171;
// bram[43508] = 150;
// bram[43509] = 128;
// bram[43510] = 107;
// bram[43511] = 85;
// bram[43512] = 65;
// bram[43513] = 47;
// bram[43514] = 31;
// bram[43515] = 18;
// bram[43516] = 8;
// bram[43517] = 2;
// bram[43518] = 0;
// bram[43519] = 1;
// bram[43520] = 6;
// bram[43521] = 14;
// bram[43522] = 26;
// bram[43523] = 41;
// bram[43524] = 58;
// bram[43525] = 78;
// bram[43526] = 99;
// bram[43527] = 121;
// bram[43528] = 142;
// bram[43529] = 164;
// bram[43530] = 184;
// bram[43531] = 203;
// bram[43532] = 219;
// bram[43533] = 233;
// bram[43534] = 243;
// bram[43535] = 250;
// bram[43536] = 253;
// bram[43537] = 253;
// bram[43538] = 248;
// bram[43539] = 241;
// bram[43540] = 229;
// bram[43541] = 215;
// bram[43542] = 198;
// bram[43543] = 179;
// bram[43544] = 158;
// bram[43545] = 136;
// bram[43546] = 115;
// bram[43547] = 93;
// bram[43548] = 72;
// bram[43549] = 53;
// bram[43550] = 37;
// bram[43551] = 23;
// bram[43552] = 12;
// bram[43553] = 4;
// bram[43554] = 0;
// bram[43555] = 0;
// bram[43556] = 3;
// bram[43557] = 11;
// bram[43558] = 21;
// bram[43559] = 35;
// bram[43560] = 52;
// bram[43561] = 71;
// bram[43562] = 91;
// bram[43563] = 113;
// bram[43564] = 134;
// bram[43565] = 156;
// bram[43566] = 177;
// bram[43567] = 196;
// bram[43568] = 213;
// bram[43569] = 228;
// bram[43570] = 240;
// bram[43571] = 248;
// bram[43572] = 252;
// bram[43573] = 253;
// bram[43574] = 250;
// bram[43575] = 244;
// bram[43576] = 234;
// bram[43577] = 220;
// bram[43578] = 204;
// bram[43579] = 186;
// bram[43580] = 166;
// bram[43581] = 144;
// bram[43582] = 123;
// bram[43583] = 101;
// bram[43584] = 80;
// bram[43585] = 60;
// bram[43586] = 43;
// bram[43587] = 27;
// bram[43588] = 15;
// bram[43589] = 6;
// bram[43590] = 1;
// bram[43591] = 0;
// bram[43592] = 2;
// bram[43593] = 8;
// bram[43594] = 17;
// bram[43595] = 30;
// bram[43596] = 46;
// bram[43597] = 64;
// bram[43598] = 83;
// bram[43599] = 105;
// bram[43600] = 127;
// bram[43601] = 148;
// bram[43602] = 170;
// bram[43603] = 189;
// bram[43604] = 207;
// bram[43605] = 223;
// bram[43606] = 236;
// bram[43607] = 245;
// bram[43608] = 251;
// bram[43609] = 253;
// bram[43610] = 252;
// bram[43611] = 247;
// bram[43612] = 238;
// bram[43613] = 226;
// bram[43614] = 210;
// bram[43615] = 193;
// bram[43616] = 173;
// bram[43617] = 152;
// bram[43618] = 130;
// bram[43619] = 109;
// bram[43620] = 87;
// bram[43621] = 67;
// bram[43622] = 49;
// bram[43623] = 33;
// bram[43624] = 19;
// bram[43625] = 9;
// bram[43626] = 3;
// bram[43627] = 0;
// bram[43628] = 1;
// bram[43629] = 5;
// bram[43630] = 13;
// bram[43631] = 25;
// bram[43632] = 40;
// bram[43633] = 57;
// bram[43634] = 76;
// bram[43635] = 97;
// bram[43636] = 119;
// bram[43637] = 140;
// bram[43638] = 162;
// bram[43639] = 182;
// bram[43640] = 201;
// bram[43641] = 218;
// bram[43642] = 232;
// bram[43643] = 242;
// bram[43644] = 250;
// bram[43645] = 253;
// bram[43646] = 253;
// bram[43647] = 249;
// bram[43648] = 241;
// bram[43649] = 230;
// bram[43650] = 216;
// bram[43651] = 200;
// bram[43652] = 181;
// bram[43653] = 160;
// bram[43654] = 138;
// bram[43655] = 117;
// bram[43656] = 95;
// bram[43657] = 74;
// bram[43658] = 55;
// bram[43659] = 38;
// bram[43660] = 24;
// bram[43661] = 12;
// bram[43662] = 5;
// bram[43663] = 0;
// bram[43664] = 0;
// bram[43665] = 3;
// bram[43666] = 10;
// bram[43667] = 20;
// bram[43668] = 34;
// bram[43669] = 50;
// bram[43670] = 69;
// bram[43671] = 89;
// bram[43672] = 111;
// bram[43673] = 132;
// bram[43674] = 154;
// bram[43675] = 175;
// bram[43676] = 195;
// bram[43677] = 212;
// bram[43678] = 227;
// bram[43679] = 239;
// bram[43680] = 247;
// bram[43681] = 252;
// bram[43682] = 253;
// bram[43683] = 251;
// bram[43684] = 245;
// bram[43685] = 235;
// bram[43686] = 222;
// bram[43687] = 206;
// bram[43688] = 188;
// bram[43689] = 168;
// bram[43690] = 146;
// bram[43691] = 125;
// bram[43692] = 103;
// bram[43693] = 82;
// bram[43694] = 62;
// bram[43695] = 44;
// bram[43696] = 29;
// bram[43697] = 16;
// bram[43698] = 7;
// bram[43699] = 1;
// bram[43700] = 0;
// bram[43701] = 1;
// bram[43702] = 7;
// bram[43703] = 16;
// bram[43704] = 29;
// bram[43705] = 44;
// bram[43706] = 62;
// bram[43707] = 82;
// bram[43708] = 103;
// bram[43709] = 125;
// bram[43710] = 146;
// bram[43711] = 168;
// bram[43712] = 188;
// bram[43713] = 206;
// bram[43714] = 222;
// bram[43715] = 235;
// bram[43716] = 245;
// bram[43717] = 251;
// bram[43718] = 253;
// bram[43719] = 252;
// bram[43720] = 247;
// bram[43721] = 239;
// bram[43722] = 227;
// bram[43723] = 212;
// bram[43724] = 195;
// bram[43725] = 175;
// bram[43726] = 154;
// bram[43727] = 132;
// bram[43728] = 111;
// bram[43729] = 89;
// bram[43730] = 69;
// bram[43731] = 50;
// bram[43732] = 34;
// bram[43733] = 20;
// bram[43734] = 10;
// bram[43735] = 3;
// bram[43736] = 0;
// bram[43737] = 0;
// bram[43738] = 5;
// bram[43739] = 12;
// bram[43740] = 24;
// bram[43741] = 38;
// bram[43742] = 55;
// bram[43743] = 74;
// bram[43744] = 95;
// bram[43745] = 117;
// bram[43746] = 138;
// bram[43747] = 160;
// bram[43748] = 181;
// bram[43749] = 200;
// bram[43750] = 216;
// bram[43751] = 230;
// bram[43752] = 241;
// bram[43753] = 249;
// bram[43754] = 253;
// bram[43755] = 253;
// bram[43756] = 250;
// bram[43757] = 242;
// bram[43758] = 232;
// bram[43759] = 218;
// bram[43760] = 201;
// bram[43761] = 182;
// bram[43762] = 162;
// bram[43763] = 140;
// bram[43764] = 119;
// bram[43765] = 97;
// bram[43766] = 76;
// bram[43767] = 57;
// bram[43768] = 40;
// bram[43769] = 25;
// bram[43770] = 13;
// bram[43771] = 5;
// bram[43772] = 1;
// bram[43773] = 0;
// bram[43774] = 3;
// bram[43775] = 9;
// bram[43776] = 19;
// bram[43777] = 33;
// bram[43778] = 49;
// bram[43779] = 67;
// bram[43780] = 87;
// bram[43781] = 109;
// bram[43782] = 130;
// bram[43783] = 152;
// bram[43784] = 173;
// bram[43785] = 193;
// bram[43786] = 210;
// bram[43787] = 226;
// bram[43788] = 238;
// bram[43789] = 247;
// bram[43790] = 252;
// bram[43791] = 253;
// bram[43792] = 251;
// bram[43793] = 245;
// bram[43794] = 236;
// bram[43795] = 223;
// bram[43796] = 207;
// bram[43797] = 189;
// bram[43798] = 170;
// bram[43799] = 148;
// bram[43800] = 126;
// bram[43801] = 105;
// bram[43802] = 83;
// bram[43803] = 64;
// bram[43804] = 46;
// bram[43805] = 30;
// bram[43806] = 17;
// bram[43807] = 8;
// bram[43808] = 2;
// bram[43809] = 0;
// bram[43810] = 1;
// bram[43811] = 6;
// bram[43812] = 15;
// bram[43813] = 27;
// bram[43814] = 43;
// bram[43815] = 60;
// bram[43816] = 80;
// bram[43817] = 101;
// bram[43818] = 123;
// bram[43819] = 144;
// bram[43820] = 166;
// bram[43821] = 186;
// bram[43822] = 204;
// bram[43823] = 220;
// bram[43824] = 234;
// bram[43825] = 244;
// bram[43826] = 250;
// bram[43827] = 253;
// bram[43828] = 252;
// bram[43829] = 248;
// bram[43830] = 240;
// bram[43831] = 228;
// bram[43832] = 213;
// bram[43833] = 196;
// bram[43834] = 177;
// bram[43835] = 156;
// bram[43836] = 134;
// bram[43837] = 113;
// bram[43838] = 91;
// bram[43839] = 71;
// bram[43840] = 52;
// bram[43841] = 35;
// bram[43842] = 21;
// bram[43843] = 11;
// bram[43844] = 3;
// bram[43845] = 0;
// bram[43846] = 0;
// bram[43847] = 4;
// bram[43848] = 12;
// bram[43849] = 23;
// bram[43850] = 37;
// bram[43851] = 53;
// bram[43852] = 72;
// bram[43853] = 93;
// bram[43854] = 115;
// bram[43855] = 136;
// bram[43856] = 158;
// bram[43857] = 179;
// bram[43858] = 198;
// bram[43859] = 215;
// bram[43860] = 229;
// bram[43861] = 241;
// bram[43862] = 248;
// bram[43863] = 253;
// bram[43864] = 253;
// bram[43865] = 250;
// bram[43866] = 243;
// bram[43867] = 233;
// bram[43868] = 219;
// bram[43869] = 203;
// bram[43870] = 184;
// bram[43871] = 164;
// bram[43872] = 142;
// bram[43873] = 121;
// bram[43874] = 99;
// bram[43875] = 78;
// bram[43876] = 58;
// bram[43877] = 41;
// bram[43878] = 26;
// bram[43879] = 14;
// bram[43880] = 6;
// bram[43881] = 1;
// bram[43882] = 0;
// bram[43883] = 2;
// bram[43884] = 8;
// bram[43885] = 18;
// bram[43886] = 31;
// bram[43887] = 47;
// bram[43888] = 65;
// bram[43889] = 85;
// bram[43890] = 107;
// bram[43891] = 128;
// bram[43892] = 150;
// bram[43893] = 171;
// bram[43894] = 191;
// bram[43895] = 209;
// bram[43896] = 224;
// bram[43897] = 237;
// bram[43898] = 246;
// bram[43899] = 252;
// bram[43900] = 254;
// bram[43901] = 252;
// bram[43902] = 246;
// bram[43903] = 237;
// bram[43904] = 224;
// bram[43905] = 209;
// bram[43906] = 191;
// bram[43907] = 171;
// bram[43908] = 150;
// bram[43909] = 128;
// bram[43910] = 107;
// bram[43911] = 85;
// bram[43912] = 65;
// bram[43913] = 47;
// bram[43914] = 31;
// bram[43915] = 18;
// bram[43916] = 8;
// bram[43917] = 2;
// bram[43918] = 0;
// bram[43919] = 1;
// bram[43920] = 6;
// bram[43921] = 14;
// bram[43922] = 26;
// bram[43923] = 41;
// bram[43924] = 58;
// bram[43925] = 78;
// bram[43926] = 99;
// bram[43927] = 121;
// bram[43928] = 142;
// bram[43929] = 164;
// bram[43930] = 184;
// bram[43931] = 203;
// bram[43932] = 219;
// bram[43933] = 233;
// bram[43934] = 243;
// bram[43935] = 250;
// bram[43936] = 253;
// bram[43937] = 253;
// bram[43938] = 248;
// bram[43939] = 241;
// bram[43940] = 229;
// bram[43941] = 215;
// bram[43942] = 198;
// bram[43943] = 179;
// bram[43944] = 158;
// bram[43945] = 136;
// bram[43946] = 115;
// bram[43947] = 93;
// bram[43948] = 72;
// bram[43949] = 53;
// bram[43950] = 37;
// bram[43951] = 23;
// bram[43952] = 12;
// bram[43953] = 4;
// bram[43954] = 0;
// bram[43955] = 0;
// bram[43956] = 3;
// bram[43957] = 11;
// bram[43958] = 21;
// bram[43959] = 35;
// bram[43960] = 52;
// bram[43961] = 71;
// bram[43962] = 91;
// bram[43963] = 113;
// bram[43964] = 134;
// bram[43965] = 156;
// bram[43966] = 177;
// bram[43967] = 196;
// bram[43968] = 213;
// bram[43969] = 228;
// bram[43970] = 240;
// bram[43971] = 248;
// bram[43972] = 252;
// bram[43973] = 253;
// bram[43974] = 250;
// bram[43975] = 244;
// bram[43976] = 234;
// bram[43977] = 220;
// bram[43978] = 204;
// bram[43979] = 186;
// bram[43980] = 166;
// bram[43981] = 144;
// bram[43982] = 123;
// bram[43983] = 101;
// bram[43984] = 80;
// bram[43985] = 60;
// bram[43986] = 43;
// bram[43987] = 27;
// bram[43988] = 15;
// bram[43989] = 6;
// bram[43990] = 1;
// bram[43991] = 0;
// bram[43992] = 2;
// bram[43993] = 8;
// bram[43994] = 17;
// bram[43995] = 30;
// bram[43996] = 46;
// bram[43997] = 64;
// bram[43998] = 83;
// bram[43999] = 105;
// bram[44000] = 127;
// bram[44001] = 148;
// bram[44002] = 170;
// bram[44003] = 189;
// bram[44004] = 207;
// bram[44005] = 223;
// bram[44006] = 236;
// bram[44007] = 245;
// bram[44008] = 251;
// bram[44009] = 253;
// bram[44010] = 252;
// bram[44011] = 247;
// bram[44012] = 238;
// bram[44013] = 226;
// bram[44014] = 210;
// bram[44015] = 193;
// bram[44016] = 173;
// bram[44017] = 152;
// bram[44018] = 130;
// bram[44019] = 109;
// bram[44020] = 87;
// bram[44021] = 67;
// bram[44022] = 49;
// bram[44023] = 33;
// bram[44024] = 19;
// bram[44025] = 9;
// bram[44026] = 3;
// bram[44027] = 0;
// bram[44028] = 1;
// bram[44029] = 5;
// bram[44030] = 13;
// bram[44031] = 25;
// bram[44032] = 40;
// bram[44033] = 57;
// bram[44034] = 76;
// bram[44035] = 97;
// bram[44036] = 119;
// bram[44037] = 140;
// bram[44038] = 162;
// bram[44039] = 182;
// bram[44040] = 201;
// bram[44041] = 218;
// bram[44042] = 232;
// bram[44043] = 242;
// bram[44044] = 250;
// bram[44045] = 253;
// bram[44046] = 253;
// bram[44047] = 249;
// bram[44048] = 241;
// bram[44049] = 230;
// bram[44050] = 216;
// bram[44051] = 200;
// bram[44052] = 181;
// bram[44053] = 160;
// bram[44054] = 138;
// bram[44055] = 117;
// bram[44056] = 95;
// bram[44057] = 74;
// bram[44058] = 55;
// bram[44059] = 38;
// bram[44060] = 24;
// bram[44061] = 12;
// bram[44062] = 5;
// bram[44063] = 0;
// bram[44064] = 0;
// bram[44065] = 3;
// bram[44066] = 10;
// bram[44067] = 20;
// bram[44068] = 34;
// bram[44069] = 50;
// bram[44070] = 69;
// bram[44071] = 89;
// bram[44072] = 111;
// bram[44073] = 132;
// bram[44074] = 154;
// bram[44075] = 175;
// bram[44076] = 195;
// bram[44077] = 212;
// bram[44078] = 227;
// bram[44079] = 239;
// bram[44080] = 247;
// bram[44081] = 252;
// bram[44082] = 253;
// bram[44083] = 251;
// bram[44084] = 245;
// bram[44085] = 235;
// bram[44086] = 222;
// bram[44087] = 206;
// bram[44088] = 188;
// bram[44089] = 168;
// bram[44090] = 146;
// bram[44091] = 125;
// bram[44092] = 103;
// bram[44093] = 82;
// bram[44094] = 62;
// bram[44095] = 44;
// bram[44096] = 29;
// bram[44097] = 16;
// bram[44098] = 7;
// bram[44099] = 1;
// bram[44100] = 0;
// bram[44101] = 1;
// bram[44102] = 7;
// bram[44103] = 16;
// bram[44104] = 29;
// bram[44105] = 44;
// bram[44106] = 62;
// bram[44107] = 82;
// bram[44108] = 103;
// bram[44109] = 125;
// bram[44110] = 146;
// bram[44111] = 168;
// bram[44112] = 188;
// bram[44113] = 206;
// bram[44114] = 222;
// bram[44115] = 235;
// bram[44116] = 245;
// bram[44117] = 251;
// bram[44118] = 253;
// bram[44119] = 252;
// bram[44120] = 247;
// bram[44121] = 239;
// bram[44122] = 227;
// bram[44123] = 212;
// bram[44124] = 195;
// bram[44125] = 175;
// bram[44126] = 154;
// bram[44127] = 132;
// bram[44128] = 111;
// bram[44129] = 89;
// bram[44130] = 69;
// bram[44131] = 50;
// bram[44132] = 34;
// bram[44133] = 20;
// bram[44134] = 10;
// bram[44135] = 3;
// bram[44136] = 0;
// bram[44137] = 0;
// bram[44138] = 5;
// bram[44139] = 12;
// bram[44140] = 24;
// bram[44141] = 38;
// bram[44142] = 55;
// bram[44143] = 74;
// bram[44144] = 95;
// bram[44145] = 117;
// bram[44146] = 138;
// bram[44147] = 160;
// bram[44148] = 181;
// bram[44149] = 200;
// bram[44150] = 216;
// bram[44151] = 230;
// bram[44152] = 241;
// bram[44153] = 249;
// bram[44154] = 253;
// bram[44155] = 253;
// bram[44156] = 250;
// bram[44157] = 242;
// bram[44158] = 232;
// bram[44159] = 218;
// bram[44160] = 201;
// bram[44161] = 182;
// bram[44162] = 162;
// bram[44163] = 140;
// bram[44164] = 119;
// bram[44165] = 97;
// bram[44166] = 76;
// bram[44167] = 57;
// bram[44168] = 40;
// bram[44169] = 25;
// bram[44170] = 13;
// bram[44171] = 5;
// bram[44172] = 1;
// bram[44173] = 0;
// bram[44174] = 3;
// bram[44175] = 9;
// bram[44176] = 19;
// bram[44177] = 33;
// bram[44178] = 49;
// bram[44179] = 67;
// bram[44180] = 87;
// bram[44181] = 109;
// bram[44182] = 130;
// bram[44183] = 152;
// bram[44184] = 173;
// bram[44185] = 193;
// bram[44186] = 210;
// bram[44187] = 226;
// bram[44188] = 238;
// bram[44189] = 247;
// bram[44190] = 252;
// bram[44191] = 253;
// bram[44192] = 251;
// bram[44193] = 245;
// bram[44194] = 236;
// bram[44195] = 223;
// bram[44196] = 207;
// bram[44197] = 189;
// bram[44198] = 170;
// bram[44199] = 148;
// bram[44200] = 126;
// bram[44201] = 105;
// bram[44202] = 83;
// bram[44203] = 64;
// bram[44204] = 46;
// bram[44205] = 30;
// bram[44206] = 17;
// bram[44207] = 8;
// bram[44208] = 2;
// bram[44209] = 0;
// bram[44210] = 1;
// bram[44211] = 6;
// bram[44212] = 15;
// bram[44213] = 27;
// bram[44214] = 43;
// bram[44215] = 60;
// bram[44216] = 80;
// bram[44217] = 101;
// bram[44218] = 123;
// bram[44219] = 144;
// bram[44220] = 166;
// bram[44221] = 186;
// bram[44222] = 204;
// bram[44223] = 220;
// bram[44224] = 234;
// bram[44225] = 244;
// bram[44226] = 250;
// bram[44227] = 253;
// bram[44228] = 252;
// bram[44229] = 248;
// bram[44230] = 240;
// bram[44231] = 228;
// bram[44232] = 213;
// bram[44233] = 196;
// bram[44234] = 177;
// bram[44235] = 156;
// bram[44236] = 134;
// bram[44237] = 113;
// bram[44238] = 91;
// bram[44239] = 71;
// bram[44240] = 52;
// bram[44241] = 35;
// bram[44242] = 21;
// bram[44243] = 11;
// bram[44244] = 3;
// bram[44245] = 0;
// bram[44246] = 0;
// bram[44247] = 4;
// bram[44248] = 12;
// bram[44249] = 23;
// bram[44250] = 37;
// bram[44251] = 53;
// bram[44252] = 72;
// bram[44253] = 93;
// bram[44254] = 115;
// bram[44255] = 136;
// bram[44256] = 158;
// bram[44257] = 179;
// bram[44258] = 198;
// bram[44259] = 215;
// bram[44260] = 229;
// bram[44261] = 241;
// bram[44262] = 248;
// bram[44263] = 253;
// bram[44264] = 253;
// bram[44265] = 250;
// bram[44266] = 243;
// bram[44267] = 233;
// bram[44268] = 219;
// bram[44269] = 203;
// bram[44270] = 184;
// bram[44271] = 164;
// bram[44272] = 142;
// bram[44273] = 121;
// bram[44274] = 99;
// bram[44275] = 78;
// bram[44276] = 58;
// bram[44277] = 41;
// bram[44278] = 26;
// bram[44279] = 14;
// bram[44280] = 6;
// bram[44281] = 1;
// bram[44282] = 0;
// bram[44283] = 2;
// bram[44284] = 8;
// bram[44285] = 18;
// bram[44286] = 31;
// bram[44287] = 47;
// bram[44288] = 65;
// bram[44289] = 85;
// bram[44290] = 107;
// bram[44291] = 128;
// bram[44292] = 150;
// bram[44293] = 171;
// bram[44294] = 191;
// bram[44295] = 209;
// bram[44296] = 224;
// bram[44297] = 237;
// bram[44298] = 246;
// bram[44299] = 252;
// bram[44300] = 254;
// bram[44301] = 252;
// bram[44302] = 246;
// bram[44303] = 237;
// bram[44304] = 224;
// bram[44305] = 209;
// bram[44306] = 191;
// bram[44307] = 171;
// bram[44308] = 150;
// bram[44309] = 128;
// bram[44310] = 107;
// bram[44311] = 85;
// bram[44312] = 65;
// bram[44313] = 47;
// bram[44314] = 31;
// bram[44315] = 18;
// bram[44316] = 8;
// bram[44317] = 2;
// bram[44318] = 0;
// bram[44319] = 1;
// bram[44320] = 6;
// bram[44321] = 14;
// bram[44322] = 26;
// bram[44323] = 41;
// bram[44324] = 58;
// bram[44325] = 78;
// bram[44326] = 99;
// bram[44327] = 121;
// bram[44328] = 142;
// bram[44329] = 164;
// bram[44330] = 184;
// bram[44331] = 203;
// bram[44332] = 219;
// bram[44333] = 233;
// bram[44334] = 243;
// bram[44335] = 250;
// bram[44336] = 253;
// bram[44337] = 253;
// bram[44338] = 248;
// bram[44339] = 241;
// bram[44340] = 229;
// bram[44341] = 215;
// bram[44342] = 198;
// bram[44343] = 179;
// bram[44344] = 158;
// bram[44345] = 136;
// bram[44346] = 115;
// bram[44347] = 93;
// bram[44348] = 72;
// bram[44349] = 53;
// bram[44350] = 37;
// bram[44351] = 23;
// bram[44352] = 12;
// bram[44353] = 4;
// bram[44354] = 0;
// bram[44355] = 0;
// bram[44356] = 3;
// bram[44357] = 11;
// bram[44358] = 21;
// bram[44359] = 35;
// bram[44360] = 52;
// bram[44361] = 71;
// bram[44362] = 91;
// bram[44363] = 113;
// bram[44364] = 134;
// bram[44365] = 156;
// bram[44366] = 177;
// bram[44367] = 196;
// bram[44368] = 213;
// bram[44369] = 228;
// bram[44370] = 240;
// bram[44371] = 248;
// bram[44372] = 252;
// bram[44373] = 253;
// bram[44374] = 250;
// bram[44375] = 244;
// bram[44376] = 234;
// bram[44377] = 220;
// bram[44378] = 204;
// bram[44379] = 186;
// bram[44380] = 166;
// bram[44381] = 144;
// bram[44382] = 123;
// bram[44383] = 101;
// bram[44384] = 80;
// bram[44385] = 60;
// bram[44386] = 43;
// bram[44387] = 27;
// bram[44388] = 15;
// bram[44389] = 6;
// bram[44390] = 1;
// bram[44391] = 0;
// bram[44392] = 2;
// bram[44393] = 8;
// bram[44394] = 17;
// bram[44395] = 30;
// bram[44396] = 46;
// bram[44397] = 64;
// bram[44398] = 83;
// bram[44399] = 105;
// bram[44400] = 127;
// bram[44401] = 148;
// bram[44402] = 170;
// bram[44403] = 189;
// bram[44404] = 207;
// bram[44405] = 223;
// bram[44406] = 236;
// bram[44407] = 245;
// bram[44408] = 251;
// bram[44409] = 253;
// bram[44410] = 252;
// bram[44411] = 247;
// bram[44412] = 238;
// bram[44413] = 226;
// bram[44414] = 210;
// bram[44415] = 193;
// bram[44416] = 173;
// bram[44417] = 152;
// bram[44418] = 130;
// bram[44419] = 109;
// bram[44420] = 87;
// bram[44421] = 67;
// bram[44422] = 49;
// bram[44423] = 33;
// bram[44424] = 19;
// bram[44425] = 9;
// bram[44426] = 3;
// bram[44427] = 0;
// bram[44428] = 1;
// bram[44429] = 5;
// bram[44430] = 13;
// bram[44431] = 25;
// bram[44432] = 40;
// bram[44433] = 57;
// bram[44434] = 76;
// bram[44435] = 97;
// bram[44436] = 119;
// bram[44437] = 140;
// bram[44438] = 162;
// bram[44439] = 182;
// bram[44440] = 201;
// bram[44441] = 218;
// bram[44442] = 232;
// bram[44443] = 242;
// bram[44444] = 250;
// bram[44445] = 253;
// bram[44446] = 253;
// bram[44447] = 249;
// bram[44448] = 241;
// bram[44449] = 230;
// bram[44450] = 216;
// bram[44451] = 200;
// bram[44452] = 181;
// bram[44453] = 160;
// bram[44454] = 138;
// bram[44455] = 117;
// bram[44456] = 95;
// bram[44457] = 74;
// bram[44458] = 55;
// bram[44459] = 38;
// bram[44460] = 24;
// bram[44461] = 12;
// bram[44462] = 5;
// bram[44463] = 0;
// bram[44464] = 0;
// bram[44465] = 3;
// bram[44466] = 10;
// bram[44467] = 20;
// bram[44468] = 34;
// bram[44469] = 50;
// bram[44470] = 69;
// bram[44471] = 89;
// bram[44472] = 111;
// bram[44473] = 132;
// bram[44474] = 154;
// bram[44475] = 175;
// bram[44476] = 195;
// bram[44477] = 212;
// bram[44478] = 227;
// bram[44479] = 239;
// bram[44480] = 247;
// bram[44481] = 252;
// bram[44482] = 253;
// bram[44483] = 251;
// bram[44484] = 245;
// bram[44485] = 235;
// bram[44486] = 222;
// bram[44487] = 206;
// bram[44488] = 188;
// bram[44489] = 168;
// bram[44490] = 146;
// bram[44491] = 125;
// bram[44492] = 103;
// bram[44493] = 82;
// bram[44494] = 62;
// bram[44495] = 44;
// bram[44496] = 29;
// bram[44497] = 16;
// bram[44498] = 7;
// bram[44499] = 1;
// bram[44500] = 0;
// bram[44501] = 1;
// bram[44502] = 7;
// bram[44503] = 16;
// bram[44504] = 29;
// bram[44505] = 44;
// bram[44506] = 62;
// bram[44507] = 82;
// bram[44508] = 103;
// bram[44509] = 125;
// bram[44510] = 146;
// bram[44511] = 168;
// bram[44512] = 188;
// bram[44513] = 206;
// bram[44514] = 222;
// bram[44515] = 235;
// bram[44516] = 245;
// bram[44517] = 251;
// bram[44518] = 253;
// bram[44519] = 252;
// bram[44520] = 247;
// bram[44521] = 239;
// bram[44522] = 227;
// bram[44523] = 212;
// bram[44524] = 195;
// bram[44525] = 175;
// bram[44526] = 154;
// bram[44527] = 132;
// bram[44528] = 111;
// bram[44529] = 89;
// bram[44530] = 69;
// bram[44531] = 50;
// bram[44532] = 34;
// bram[44533] = 20;
// bram[44534] = 10;
// bram[44535] = 3;
// bram[44536] = 0;
// bram[44537] = 0;
// bram[44538] = 5;
// bram[44539] = 12;
// bram[44540] = 24;
// bram[44541] = 38;
// bram[44542] = 55;
// bram[44543] = 74;
// bram[44544] = 95;
// bram[44545] = 117;
// bram[44546] = 138;
// bram[44547] = 160;
// bram[44548] = 181;
// bram[44549] = 200;
// bram[44550] = 216;
// bram[44551] = 230;
// bram[44552] = 241;
// bram[44553] = 249;
// bram[44554] = 253;
// bram[44555] = 253;
// bram[44556] = 250;
// bram[44557] = 242;
// bram[44558] = 232;
// bram[44559] = 218;
// bram[44560] = 201;
// bram[44561] = 182;
// bram[44562] = 162;
// bram[44563] = 140;
// bram[44564] = 119;
// bram[44565] = 97;
// bram[44566] = 76;
// bram[44567] = 57;
// bram[44568] = 40;
// bram[44569] = 25;
// bram[44570] = 13;
// bram[44571] = 5;
// bram[44572] = 1;
// bram[44573] = 0;
// bram[44574] = 3;
// bram[44575] = 9;
// bram[44576] = 19;
// bram[44577] = 33;
// bram[44578] = 49;
// bram[44579] = 67;
// bram[44580] = 87;
// bram[44581] = 109;
// bram[44582] = 130;
// bram[44583] = 152;
// bram[44584] = 173;
// bram[44585] = 193;
// bram[44586] = 210;
// bram[44587] = 226;
// bram[44588] = 238;
// bram[44589] = 247;
// bram[44590] = 252;
// bram[44591] = 253;
// bram[44592] = 251;
// bram[44593] = 245;
// bram[44594] = 236;
// bram[44595] = 223;
// bram[44596] = 207;
// bram[44597] = 189;
// bram[44598] = 170;
// bram[44599] = 148;
// bram[44600] = 126;
// bram[44601] = 105;
// bram[44602] = 83;
// bram[44603] = 64;
// bram[44604] = 46;
// bram[44605] = 30;
// bram[44606] = 17;
// bram[44607] = 8;
// bram[44608] = 2;
// bram[44609] = 0;
// bram[44610] = 1;
// bram[44611] = 6;
// bram[44612] = 15;
// bram[44613] = 27;
// bram[44614] = 43;
// bram[44615] = 60;
// bram[44616] = 80;
// bram[44617] = 101;
// bram[44618] = 123;
// bram[44619] = 144;
// bram[44620] = 166;
// bram[44621] = 186;
// bram[44622] = 204;
// bram[44623] = 220;
// bram[44624] = 234;
// bram[44625] = 244;
// bram[44626] = 250;
// bram[44627] = 253;
// bram[44628] = 252;
// bram[44629] = 248;
// bram[44630] = 240;
// bram[44631] = 228;
// bram[44632] = 213;
// bram[44633] = 196;
// bram[44634] = 177;
// bram[44635] = 156;
// bram[44636] = 134;
// bram[44637] = 113;
// bram[44638] = 91;
// bram[44639] = 71;
// bram[44640] = 52;
// bram[44641] = 35;
// bram[44642] = 21;
// bram[44643] = 11;
// bram[44644] = 3;
// bram[44645] = 0;
// bram[44646] = 0;
// bram[44647] = 4;
// bram[44648] = 12;
// bram[44649] = 23;
// bram[44650] = 37;
// bram[44651] = 53;
// bram[44652] = 72;
// bram[44653] = 93;
// bram[44654] = 115;
// bram[44655] = 136;
// bram[44656] = 158;
// bram[44657] = 179;
// bram[44658] = 198;
// bram[44659] = 215;
// bram[44660] = 229;
// bram[44661] = 241;
// bram[44662] = 248;
// bram[44663] = 253;
// bram[44664] = 253;
// bram[44665] = 250;
// bram[44666] = 243;
// bram[44667] = 233;
// bram[44668] = 219;
// bram[44669] = 203;
// bram[44670] = 184;
// bram[44671] = 164;
// bram[44672] = 142;
// bram[44673] = 121;
// bram[44674] = 99;
// bram[44675] = 78;
// bram[44676] = 58;
// bram[44677] = 41;
// bram[44678] = 26;
// bram[44679] = 14;
// bram[44680] = 6;
// bram[44681] = 1;
// bram[44682] = 0;
// bram[44683] = 2;
// bram[44684] = 8;
// bram[44685] = 18;
// bram[44686] = 31;
// bram[44687] = 47;
// bram[44688] = 65;
// bram[44689] = 85;
// bram[44690] = 107;
// bram[44691] = 128;
// bram[44692] = 150;
// bram[44693] = 171;
// bram[44694] = 191;
// bram[44695] = 209;
// bram[44696] = 224;
// bram[44697] = 237;
// bram[44698] = 246;
// bram[44699] = 252;
// bram[44700] = 254;
// bram[44701] = 252;
// bram[44702] = 246;
// bram[44703] = 237;
// bram[44704] = 224;
// bram[44705] = 209;
// bram[44706] = 191;
// bram[44707] = 171;
// bram[44708] = 150;
// bram[44709] = 128;
// bram[44710] = 107;
// bram[44711] = 85;
// bram[44712] = 65;
// bram[44713] = 47;
// bram[44714] = 31;
// bram[44715] = 18;
// bram[44716] = 8;
// bram[44717] = 2;
// bram[44718] = 0;
// bram[44719] = 1;
// bram[44720] = 6;
// bram[44721] = 14;
// bram[44722] = 26;
// bram[44723] = 41;
// bram[44724] = 58;
// bram[44725] = 78;
// bram[44726] = 99;
// bram[44727] = 121;
// bram[44728] = 142;
// bram[44729] = 164;
// bram[44730] = 184;
// bram[44731] = 203;
// bram[44732] = 219;
// bram[44733] = 233;
// bram[44734] = 243;
// bram[44735] = 250;
// bram[44736] = 253;
// bram[44737] = 253;
// bram[44738] = 248;
// bram[44739] = 241;
// bram[44740] = 229;
// bram[44741] = 215;
// bram[44742] = 198;
// bram[44743] = 179;
// bram[44744] = 158;
// bram[44745] = 136;
// bram[44746] = 115;
// bram[44747] = 93;
// bram[44748] = 72;
// bram[44749] = 53;
// bram[44750] = 37;
// bram[44751] = 23;
// bram[44752] = 12;
// bram[44753] = 4;
// bram[44754] = 0;
// bram[44755] = 0;
// bram[44756] = 3;
// bram[44757] = 11;
// bram[44758] = 21;
// bram[44759] = 35;
// bram[44760] = 52;
// bram[44761] = 71;
// bram[44762] = 91;
// bram[44763] = 113;
// bram[44764] = 134;
// bram[44765] = 156;
// bram[44766] = 177;
// bram[44767] = 196;
// bram[44768] = 213;
// bram[44769] = 228;
// bram[44770] = 240;
// bram[44771] = 248;
// bram[44772] = 252;
// bram[44773] = 253;
// bram[44774] = 250;
// bram[44775] = 244;
// bram[44776] = 234;
// bram[44777] = 220;
// bram[44778] = 204;
// bram[44779] = 186;
// bram[44780] = 166;
// bram[44781] = 144;
// bram[44782] = 123;
// bram[44783] = 101;
// bram[44784] = 80;
// bram[44785] = 60;
// bram[44786] = 43;
// bram[44787] = 27;
// bram[44788] = 15;
// bram[44789] = 6;
// bram[44790] = 1;
// bram[44791] = 0;
// bram[44792] = 2;
// bram[44793] = 8;
// bram[44794] = 17;
// bram[44795] = 30;
// bram[44796] = 46;
// bram[44797] = 64;
// bram[44798] = 83;
// bram[44799] = 105;
// bram[44800] = 126;
// bram[44801] = 148;
// bram[44802] = 170;
// bram[44803] = 189;
// bram[44804] = 207;
// bram[44805] = 223;
// bram[44806] = 236;
// bram[44807] = 245;
// bram[44808] = 251;
// bram[44809] = 253;
// bram[44810] = 252;
// bram[44811] = 247;
// bram[44812] = 238;
// bram[44813] = 226;
// bram[44814] = 210;
// bram[44815] = 193;
// bram[44816] = 173;
// bram[44817] = 152;
// bram[44818] = 130;
// bram[44819] = 109;
// bram[44820] = 87;
// bram[44821] = 67;
// bram[44822] = 49;
// bram[44823] = 33;
// bram[44824] = 19;
// bram[44825] = 9;
// bram[44826] = 3;
// bram[44827] = 0;
// bram[44828] = 1;
// bram[44829] = 5;
// bram[44830] = 13;
// bram[44831] = 25;
// bram[44832] = 40;
// bram[44833] = 57;
// bram[44834] = 76;
// bram[44835] = 97;
// bram[44836] = 119;
// bram[44837] = 140;
// bram[44838] = 162;
// bram[44839] = 182;
// bram[44840] = 201;
// bram[44841] = 218;
// bram[44842] = 232;
// bram[44843] = 242;
// bram[44844] = 250;
// bram[44845] = 253;
// bram[44846] = 253;
// bram[44847] = 249;
// bram[44848] = 241;
// bram[44849] = 230;
// bram[44850] = 216;
// bram[44851] = 200;
// bram[44852] = 181;
// bram[44853] = 160;
// bram[44854] = 138;
// bram[44855] = 117;
// bram[44856] = 95;
// bram[44857] = 74;
// bram[44858] = 55;
// bram[44859] = 38;
// bram[44860] = 24;
// bram[44861] = 12;
// bram[44862] = 5;
// bram[44863] = 0;
// bram[44864] = 0;
// bram[44865] = 3;
// bram[44866] = 10;
// bram[44867] = 20;
// bram[44868] = 34;
// bram[44869] = 50;
// bram[44870] = 69;
// bram[44871] = 89;
// bram[44872] = 111;
// bram[44873] = 132;
// bram[44874] = 154;
// bram[44875] = 175;
// bram[44876] = 195;
// bram[44877] = 212;
// bram[44878] = 227;
// bram[44879] = 239;
// bram[44880] = 247;
// bram[44881] = 252;
// bram[44882] = 253;
// bram[44883] = 251;
// bram[44884] = 245;
// bram[44885] = 235;
// bram[44886] = 222;
// bram[44887] = 206;
// bram[44888] = 188;
// bram[44889] = 168;
// bram[44890] = 146;
// bram[44891] = 125;
// bram[44892] = 103;
// bram[44893] = 82;
// bram[44894] = 62;
// bram[44895] = 44;
// bram[44896] = 29;
// bram[44897] = 16;
// bram[44898] = 7;
// bram[44899] = 1;
// bram[44900] = 0;
// bram[44901] = 1;
// bram[44902] = 7;
// bram[44903] = 16;
// bram[44904] = 29;
// bram[44905] = 44;
// bram[44906] = 62;
// bram[44907] = 82;
// bram[44908] = 103;
// bram[44909] = 125;
// bram[44910] = 146;
// bram[44911] = 168;
// bram[44912] = 188;
// bram[44913] = 206;
// bram[44914] = 222;
// bram[44915] = 235;
// bram[44916] = 245;
// bram[44917] = 251;
// bram[44918] = 253;
// bram[44919] = 252;
// bram[44920] = 247;
// bram[44921] = 239;
// bram[44922] = 227;
// bram[44923] = 212;
// bram[44924] = 195;
// bram[44925] = 175;
// bram[44926] = 154;
// bram[44927] = 132;
// bram[44928] = 111;
// bram[44929] = 89;
// bram[44930] = 69;
// bram[44931] = 50;
// bram[44932] = 34;
// bram[44933] = 20;
// bram[44934] = 10;
// bram[44935] = 3;
// bram[44936] = 0;
// bram[44937] = 0;
// bram[44938] = 5;
// bram[44939] = 12;
// bram[44940] = 24;
// bram[44941] = 38;
// bram[44942] = 55;
// bram[44943] = 74;
// bram[44944] = 95;
// bram[44945] = 117;
// bram[44946] = 138;
// bram[44947] = 160;
// bram[44948] = 181;
// bram[44949] = 200;
// bram[44950] = 216;
// bram[44951] = 230;
// bram[44952] = 241;
// bram[44953] = 249;
// bram[44954] = 253;
// bram[44955] = 253;
// bram[44956] = 250;
// bram[44957] = 242;
// bram[44958] = 232;
// bram[44959] = 218;
// bram[44960] = 201;
// bram[44961] = 182;
// bram[44962] = 162;
// bram[44963] = 140;
// bram[44964] = 119;
// bram[44965] = 97;
// bram[44966] = 76;
// bram[44967] = 57;
// bram[44968] = 40;
// bram[44969] = 25;
// bram[44970] = 13;
// bram[44971] = 5;
// bram[44972] = 1;
// bram[44973] = 0;
// bram[44974] = 3;
// bram[44975] = 9;
// bram[44976] = 19;
// bram[44977] = 33;
// bram[44978] = 49;
// bram[44979] = 67;
// bram[44980] = 87;
// bram[44981] = 109;
// bram[44982] = 130;
// bram[44983] = 152;
// bram[44984] = 173;
// bram[44985] = 193;
// bram[44986] = 210;
// bram[44987] = 226;
// bram[44988] = 238;
// bram[44989] = 247;
// bram[44990] = 252;
// bram[44991] = 253;
// bram[44992] = 251;
// bram[44993] = 245;
// bram[44994] = 236;
// bram[44995] = 223;
// bram[44996] = 207;
// bram[44997] = 189;
// bram[44998] = 170;
// bram[44999] = 148;
// bram[45000] = 127;
// bram[45001] = 105;
// bram[45002] = 83;
// bram[45003] = 64;
// bram[45004] = 46;
// bram[45005] = 30;
// bram[45006] = 17;
// bram[45007] = 8;
// bram[45008] = 2;
// bram[45009] = 0;
// bram[45010] = 1;
// bram[45011] = 6;
// bram[45012] = 15;
// bram[45013] = 27;
// bram[45014] = 43;
// bram[45015] = 60;
// bram[45016] = 80;
// bram[45017] = 101;
// bram[45018] = 123;
// bram[45019] = 144;
// bram[45020] = 166;
// bram[45021] = 186;
// bram[45022] = 204;
// bram[45023] = 220;
// bram[45024] = 234;
// bram[45025] = 244;
// bram[45026] = 250;
// bram[45027] = 253;
// bram[45028] = 252;
// bram[45029] = 248;
// bram[45030] = 240;
// bram[45031] = 228;
// bram[45032] = 213;
// bram[45033] = 196;
// bram[45034] = 177;
// bram[45035] = 156;
// bram[45036] = 134;
// bram[45037] = 113;
// bram[45038] = 91;
// bram[45039] = 71;
// bram[45040] = 52;
// bram[45041] = 35;
// bram[45042] = 21;
// bram[45043] = 11;
// bram[45044] = 3;
// bram[45045] = 0;
// bram[45046] = 0;
// bram[45047] = 4;
// bram[45048] = 12;
// bram[45049] = 23;
// bram[45050] = 37;
// bram[45051] = 53;
// bram[45052] = 72;
// bram[45053] = 93;
// bram[45054] = 115;
// bram[45055] = 136;
// bram[45056] = 158;
// bram[45057] = 179;
// bram[45058] = 198;
// bram[45059] = 215;
// bram[45060] = 229;
// bram[45061] = 241;
// bram[45062] = 248;
// bram[45063] = 253;
// bram[45064] = 253;
// bram[45065] = 250;
// bram[45066] = 243;
// bram[45067] = 233;
// bram[45068] = 219;
// bram[45069] = 203;
// bram[45070] = 184;
// bram[45071] = 164;
// bram[45072] = 142;
// bram[45073] = 121;
// bram[45074] = 99;
// bram[45075] = 78;
// bram[45076] = 58;
// bram[45077] = 41;
// bram[45078] = 26;
// bram[45079] = 14;
// bram[45080] = 6;
// bram[45081] = 1;
// bram[45082] = 0;
// bram[45083] = 2;
// bram[45084] = 8;
// bram[45085] = 18;
// bram[45086] = 31;
// bram[45087] = 47;
// bram[45088] = 65;
// bram[45089] = 85;
// bram[45090] = 107;
// bram[45091] = 128;
// bram[45092] = 150;
// bram[45093] = 171;
// bram[45094] = 191;
// bram[45095] = 209;
// bram[45096] = 224;
// bram[45097] = 237;
// bram[45098] = 246;
// bram[45099] = 252;
// bram[45100] = 254;
// bram[45101] = 252;
// bram[45102] = 246;
// bram[45103] = 237;
// bram[45104] = 224;
// bram[45105] = 209;
// bram[45106] = 191;
// bram[45107] = 171;
// bram[45108] = 150;
// bram[45109] = 128;
// bram[45110] = 107;
// bram[45111] = 85;
// bram[45112] = 65;
// bram[45113] = 47;
// bram[45114] = 31;
// bram[45115] = 18;
// bram[45116] = 8;
// bram[45117] = 2;
// bram[45118] = 0;
// bram[45119] = 1;
// bram[45120] = 6;
// bram[45121] = 14;
// bram[45122] = 26;
// bram[45123] = 41;
// bram[45124] = 58;
// bram[45125] = 78;
// bram[45126] = 99;
// bram[45127] = 121;
// bram[45128] = 142;
// bram[45129] = 164;
// bram[45130] = 184;
// bram[45131] = 203;
// bram[45132] = 219;
// bram[45133] = 233;
// bram[45134] = 243;
// bram[45135] = 250;
// bram[45136] = 253;
// bram[45137] = 253;
// bram[45138] = 248;
// bram[45139] = 241;
// bram[45140] = 229;
// bram[45141] = 215;
// bram[45142] = 198;
// bram[45143] = 179;
// bram[45144] = 158;
// bram[45145] = 136;
// bram[45146] = 115;
// bram[45147] = 93;
// bram[45148] = 72;
// bram[45149] = 53;
// bram[45150] = 37;
// bram[45151] = 23;
// bram[45152] = 12;
// bram[45153] = 4;
// bram[45154] = 0;
// bram[45155] = 0;
// bram[45156] = 3;
// bram[45157] = 11;
// bram[45158] = 21;
// bram[45159] = 35;
// bram[45160] = 52;
// bram[45161] = 71;
// bram[45162] = 91;
// bram[45163] = 113;
// bram[45164] = 134;
// bram[45165] = 156;
// bram[45166] = 177;
// bram[45167] = 196;
// bram[45168] = 213;
// bram[45169] = 228;
// bram[45170] = 240;
// bram[45171] = 248;
// bram[45172] = 252;
// bram[45173] = 253;
// bram[45174] = 250;
// bram[45175] = 244;
// bram[45176] = 234;
// bram[45177] = 220;
// bram[45178] = 204;
// bram[45179] = 186;
// bram[45180] = 166;
// bram[45181] = 144;
// bram[45182] = 123;
// bram[45183] = 101;
// bram[45184] = 80;
// bram[45185] = 60;
// bram[45186] = 43;
// bram[45187] = 27;
// bram[45188] = 15;
// bram[45189] = 6;
// bram[45190] = 1;
// bram[45191] = 0;
// bram[45192] = 2;
// bram[45193] = 8;
// bram[45194] = 17;
// bram[45195] = 30;
// bram[45196] = 46;
// bram[45197] = 64;
// bram[45198] = 83;
// bram[45199] = 105;
// bram[45200] = 127;
// bram[45201] = 148;
// bram[45202] = 170;
// bram[45203] = 189;
// bram[45204] = 207;
// bram[45205] = 223;
// bram[45206] = 236;
// bram[45207] = 245;
// bram[45208] = 251;
// bram[45209] = 253;
// bram[45210] = 252;
// bram[45211] = 247;
// bram[45212] = 238;
// bram[45213] = 226;
// bram[45214] = 210;
// bram[45215] = 193;
// bram[45216] = 173;
// bram[45217] = 152;
// bram[45218] = 130;
// bram[45219] = 109;
// bram[45220] = 87;
// bram[45221] = 67;
// bram[45222] = 49;
// bram[45223] = 33;
// bram[45224] = 19;
// bram[45225] = 9;
// bram[45226] = 3;
// bram[45227] = 0;
// bram[45228] = 1;
// bram[45229] = 5;
// bram[45230] = 13;
// bram[45231] = 25;
// bram[45232] = 40;
// bram[45233] = 57;
// bram[45234] = 76;
// bram[45235] = 97;
// bram[45236] = 119;
// bram[45237] = 140;
// bram[45238] = 162;
// bram[45239] = 182;
// bram[45240] = 201;
// bram[45241] = 218;
// bram[45242] = 232;
// bram[45243] = 242;
// bram[45244] = 250;
// bram[45245] = 253;
// bram[45246] = 253;
// bram[45247] = 249;
// bram[45248] = 241;
// bram[45249] = 230;
// bram[45250] = 216;
// bram[45251] = 200;
// bram[45252] = 181;
// bram[45253] = 160;
// bram[45254] = 138;
// bram[45255] = 117;
// bram[45256] = 95;
// bram[45257] = 74;
// bram[45258] = 55;
// bram[45259] = 38;
// bram[45260] = 24;
// bram[45261] = 12;
// bram[45262] = 5;
// bram[45263] = 0;
// bram[45264] = 0;
// bram[45265] = 3;
// bram[45266] = 10;
// bram[45267] = 20;
// bram[45268] = 34;
// bram[45269] = 50;
// bram[45270] = 69;
// bram[45271] = 89;
// bram[45272] = 111;
// bram[45273] = 132;
// bram[45274] = 154;
// bram[45275] = 175;
// bram[45276] = 195;
// bram[45277] = 212;
// bram[45278] = 227;
// bram[45279] = 239;
// bram[45280] = 247;
// bram[45281] = 252;
// bram[45282] = 253;
// bram[45283] = 251;
// bram[45284] = 245;
// bram[45285] = 235;
// bram[45286] = 222;
// bram[45287] = 206;
// bram[45288] = 188;
// bram[45289] = 168;
// bram[45290] = 146;
// bram[45291] = 125;
// bram[45292] = 103;
// bram[45293] = 82;
// bram[45294] = 62;
// bram[45295] = 44;
// bram[45296] = 29;
// bram[45297] = 16;
// bram[45298] = 7;
// bram[45299] = 1;
// bram[45300] = 0;
// bram[45301] = 1;
// bram[45302] = 7;
// bram[45303] = 16;
// bram[45304] = 29;
// bram[45305] = 44;
// bram[45306] = 62;
// bram[45307] = 82;
// bram[45308] = 103;
// bram[45309] = 125;
// bram[45310] = 146;
// bram[45311] = 168;
// bram[45312] = 188;
// bram[45313] = 206;
// bram[45314] = 222;
// bram[45315] = 235;
// bram[45316] = 245;
// bram[45317] = 251;
// bram[45318] = 253;
// bram[45319] = 252;
// bram[45320] = 247;
// bram[45321] = 239;
// bram[45322] = 227;
// bram[45323] = 212;
// bram[45324] = 195;
// bram[45325] = 175;
// bram[45326] = 154;
// bram[45327] = 132;
// bram[45328] = 111;
// bram[45329] = 89;
// bram[45330] = 69;
// bram[45331] = 50;
// bram[45332] = 34;
// bram[45333] = 20;
// bram[45334] = 10;
// bram[45335] = 3;
// bram[45336] = 0;
// bram[45337] = 0;
// bram[45338] = 5;
// bram[45339] = 12;
// bram[45340] = 24;
// bram[45341] = 38;
// bram[45342] = 55;
// bram[45343] = 74;
// bram[45344] = 95;
// bram[45345] = 117;
// bram[45346] = 138;
// bram[45347] = 160;
// bram[45348] = 181;
// bram[45349] = 200;
// bram[45350] = 216;
// bram[45351] = 230;
// bram[45352] = 241;
// bram[45353] = 249;
// bram[45354] = 253;
// bram[45355] = 253;
// bram[45356] = 250;
// bram[45357] = 242;
// bram[45358] = 232;
// bram[45359] = 218;
// bram[45360] = 201;
// bram[45361] = 182;
// bram[45362] = 162;
// bram[45363] = 140;
// bram[45364] = 119;
// bram[45365] = 97;
// bram[45366] = 76;
// bram[45367] = 57;
// bram[45368] = 40;
// bram[45369] = 25;
// bram[45370] = 13;
// bram[45371] = 5;
// bram[45372] = 1;
// bram[45373] = 0;
// bram[45374] = 3;
// bram[45375] = 9;
// bram[45376] = 19;
// bram[45377] = 33;
// bram[45378] = 49;
// bram[45379] = 67;
// bram[45380] = 87;
// bram[45381] = 109;
// bram[45382] = 130;
// bram[45383] = 152;
// bram[45384] = 173;
// bram[45385] = 193;
// bram[45386] = 210;
// bram[45387] = 226;
// bram[45388] = 238;
// bram[45389] = 247;
// bram[45390] = 252;
// bram[45391] = 253;
// bram[45392] = 251;
// bram[45393] = 245;
// bram[45394] = 236;
// bram[45395] = 223;
// bram[45396] = 207;
// bram[45397] = 189;
// bram[45398] = 170;
// bram[45399] = 148;
// bram[45400] = 126;
// bram[45401] = 105;
// bram[45402] = 83;
// bram[45403] = 64;
// bram[45404] = 46;
// bram[45405] = 30;
// bram[45406] = 17;
// bram[45407] = 8;
// bram[45408] = 2;
// bram[45409] = 0;
// bram[45410] = 1;
// bram[45411] = 6;
// bram[45412] = 15;
// bram[45413] = 27;
// bram[45414] = 43;
// bram[45415] = 60;
// bram[45416] = 80;
// bram[45417] = 101;
// bram[45418] = 123;
// bram[45419] = 144;
// bram[45420] = 166;
// bram[45421] = 186;
// bram[45422] = 204;
// bram[45423] = 220;
// bram[45424] = 234;
// bram[45425] = 244;
// bram[45426] = 250;
// bram[45427] = 253;
// bram[45428] = 252;
// bram[45429] = 248;
// bram[45430] = 240;
// bram[45431] = 228;
// bram[45432] = 213;
// bram[45433] = 196;
// bram[45434] = 177;
// bram[45435] = 156;
// bram[45436] = 134;
// bram[45437] = 113;
// bram[45438] = 91;
// bram[45439] = 71;
// bram[45440] = 52;
// bram[45441] = 35;
// bram[45442] = 21;
// bram[45443] = 11;
// bram[45444] = 3;
// bram[45445] = 0;
// bram[45446] = 0;
// bram[45447] = 4;
// bram[45448] = 12;
// bram[45449] = 23;
// bram[45450] = 37;
// bram[45451] = 53;
// bram[45452] = 72;
// bram[45453] = 93;
// bram[45454] = 115;
// bram[45455] = 136;
// bram[45456] = 158;
// bram[45457] = 179;
// bram[45458] = 198;
// bram[45459] = 215;
// bram[45460] = 229;
// bram[45461] = 241;
// bram[45462] = 248;
// bram[45463] = 253;
// bram[45464] = 253;
// bram[45465] = 250;
// bram[45466] = 243;
// bram[45467] = 233;
// bram[45468] = 219;
// bram[45469] = 203;
// bram[45470] = 184;
// bram[45471] = 164;
// bram[45472] = 142;
// bram[45473] = 121;
// bram[45474] = 99;
// bram[45475] = 78;
// bram[45476] = 58;
// bram[45477] = 41;
// bram[45478] = 26;
// bram[45479] = 14;
// bram[45480] = 6;
// bram[45481] = 1;
// bram[45482] = 0;
// bram[45483] = 2;
// bram[45484] = 8;
// bram[45485] = 18;
// bram[45486] = 31;
// bram[45487] = 47;
// bram[45488] = 65;
// bram[45489] = 85;
// bram[45490] = 107;
// bram[45491] = 128;
// bram[45492] = 150;
// bram[45493] = 171;
// bram[45494] = 191;
// bram[45495] = 209;
// bram[45496] = 224;
// bram[45497] = 237;
// bram[45498] = 246;
// bram[45499] = 252;
// bram[45500] = 254;
// bram[45501] = 252;
// bram[45502] = 246;
// bram[45503] = 237;
// bram[45504] = 224;
// bram[45505] = 209;
// bram[45506] = 191;
// bram[45507] = 171;
// bram[45508] = 150;
// bram[45509] = 128;
// bram[45510] = 107;
// bram[45511] = 85;
// bram[45512] = 65;
// bram[45513] = 47;
// bram[45514] = 31;
// bram[45515] = 18;
// bram[45516] = 8;
// bram[45517] = 2;
// bram[45518] = 0;
// bram[45519] = 1;
// bram[45520] = 6;
// bram[45521] = 14;
// bram[45522] = 26;
// bram[45523] = 41;
// bram[45524] = 58;
// bram[45525] = 78;
// bram[45526] = 99;
// bram[45527] = 121;
// bram[45528] = 142;
// bram[45529] = 164;
// bram[45530] = 184;
// bram[45531] = 203;
// bram[45532] = 219;
// bram[45533] = 233;
// bram[45534] = 243;
// bram[45535] = 250;
// bram[45536] = 253;
// bram[45537] = 253;
// bram[45538] = 248;
// bram[45539] = 241;
// bram[45540] = 229;
// bram[45541] = 215;
// bram[45542] = 198;
// bram[45543] = 179;
// bram[45544] = 158;
// bram[45545] = 136;
// bram[45546] = 115;
// bram[45547] = 93;
// bram[45548] = 72;
// bram[45549] = 53;
// bram[45550] = 37;
// bram[45551] = 23;
// bram[45552] = 12;
// bram[45553] = 4;
// bram[45554] = 0;
// bram[45555] = 0;
// bram[45556] = 3;
// bram[45557] = 11;
// bram[45558] = 21;
// bram[45559] = 35;
// bram[45560] = 52;
// bram[45561] = 71;
// bram[45562] = 91;
// bram[45563] = 113;
// bram[45564] = 134;
// bram[45565] = 156;
// bram[45566] = 177;
// bram[45567] = 196;
// bram[45568] = 213;
// bram[45569] = 228;
// bram[45570] = 240;
// bram[45571] = 248;
// bram[45572] = 252;
// bram[45573] = 253;
// bram[45574] = 250;
// bram[45575] = 244;
// bram[45576] = 234;
// bram[45577] = 220;
// bram[45578] = 204;
// bram[45579] = 186;
// bram[45580] = 166;
// bram[45581] = 144;
// bram[45582] = 123;
// bram[45583] = 101;
// bram[45584] = 80;
// bram[45585] = 60;
// bram[45586] = 43;
// bram[45587] = 27;
// bram[45588] = 15;
// bram[45589] = 6;
// bram[45590] = 1;
// bram[45591] = 0;
// bram[45592] = 2;
// bram[45593] = 8;
// bram[45594] = 17;
// bram[45595] = 30;
// bram[45596] = 46;
// bram[45597] = 64;
// bram[45598] = 83;
// bram[45599] = 105;
// bram[45600] = 127;
// bram[45601] = 148;
// bram[45602] = 170;
// bram[45603] = 189;
// bram[45604] = 207;
// bram[45605] = 223;
// bram[45606] = 236;
// bram[45607] = 245;
// bram[45608] = 251;
// bram[45609] = 253;
// bram[45610] = 252;
// bram[45611] = 247;
// bram[45612] = 238;
// bram[45613] = 226;
// bram[45614] = 210;
// bram[45615] = 193;
// bram[45616] = 173;
// bram[45617] = 152;
// bram[45618] = 130;
// bram[45619] = 109;
// bram[45620] = 87;
// bram[45621] = 67;
// bram[45622] = 49;
// bram[45623] = 33;
// bram[45624] = 19;
// bram[45625] = 9;
// bram[45626] = 3;
// bram[45627] = 0;
// bram[45628] = 1;
// bram[45629] = 5;
// bram[45630] = 13;
// bram[45631] = 25;
// bram[45632] = 40;
// bram[45633] = 57;
// bram[45634] = 76;
// bram[45635] = 97;
// bram[45636] = 119;
// bram[45637] = 140;
// bram[45638] = 162;
// bram[45639] = 182;
// bram[45640] = 201;
// bram[45641] = 218;
// bram[45642] = 232;
// bram[45643] = 242;
// bram[45644] = 250;
// bram[45645] = 253;
// bram[45646] = 253;
// bram[45647] = 249;
// bram[45648] = 241;
// bram[45649] = 230;
// bram[45650] = 216;
// bram[45651] = 200;
// bram[45652] = 181;
// bram[45653] = 160;
// bram[45654] = 138;
// bram[45655] = 117;
// bram[45656] = 95;
// bram[45657] = 74;
// bram[45658] = 55;
// bram[45659] = 38;
// bram[45660] = 24;
// bram[45661] = 12;
// bram[45662] = 5;
// bram[45663] = 0;
// bram[45664] = 0;
// bram[45665] = 3;
// bram[45666] = 10;
// bram[45667] = 20;
// bram[45668] = 34;
// bram[45669] = 50;
// bram[45670] = 69;
// bram[45671] = 89;
// bram[45672] = 111;
// bram[45673] = 132;
// bram[45674] = 154;
// bram[45675] = 175;
// bram[45676] = 195;
// bram[45677] = 212;
// bram[45678] = 227;
// bram[45679] = 239;
// bram[45680] = 247;
// bram[45681] = 252;
// bram[45682] = 253;
// bram[45683] = 251;
// bram[45684] = 245;
// bram[45685] = 235;
// bram[45686] = 222;
// bram[45687] = 206;
// bram[45688] = 188;
// bram[45689] = 168;
// bram[45690] = 146;
// bram[45691] = 125;
// bram[45692] = 103;
// bram[45693] = 82;
// bram[45694] = 62;
// bram[45695] = 44;
// bram[45696] = 29;
// bram[45697] = 16;
// bram[45698] = 7;
// bram[45699] = 1;
// bram[45700] = 0;
// bram[45701] = 1;
// bram[45702] = 7;
// bram[45703] = 16;
// bram[45704] = 29;
// bram[45705] = 44;
// bram[45706] = 62;
// bram[45707] = 82;
// bram[45708] = 103;
// bram[45709] = 125;
// bram[45710] = 146;
// bram[45711] = 168;
// bram[45712] = 188;
// bram[45713] = 206;
// bram[45714] = 222;
// bram[45715] = 235;
// bram[45716] = 245;
// bram[45717] = 251;
// bram[45718] = 253;
// bram[45719] = 252;
// bram[45720] = 247;
// bram[45721] = 239;
// bram[45722] = 227;
// bram[45723] = 212;
// bram[45724] = 195;
// bram[45725] = 175;
// bram[45726] = 154;
// bram[45727] = 132;
// bram[45728] = 111;
// bram[45729] = 89;
// bram[45730] = 69;
// bram[45731] = 50;
// bram[45732] = 34;
// bram[45733] = 20;
// bram[45734] = 10;
// bram[45735] = 3;
// bram[45736] = 0;
// bram[45737] = 0;
// bram[45738] = 5;
// bram[45739] = 12;
// bram[45740] = 24;
// bram[45741] = 38;
// bram[45742] = 55;
// bram[45743] = 74;
// bram[45744] = 95;
// bram[45745] = 117;
// bram[45746] = 138;
// bram[45747] = 160;
// bram[45748] = 181;
// bram[45749] = 200;
// bram[45750] = 216;
// bram[45751] = 230;
// bram[45752] = 241;
// bram[45753] = 249;
// bram[45754] = 253;
// bram[45755] = 253;
// bram[45756] = 250;
// bram[45757] = 242;
// bram[45758] = 232;
// bram[45759] = 218;
// bram[45760] = 201;
// bram[45761] = 182;
// bram[45762] = 162;
// bram[45763] = 140;
// bram[45764] = 119;
// bram[45765] = 97;
// bram[45766] = 76;
// bram[45767] = 57;
// bram[45768] = 40;
// bram[45769] = 25;
// bram[45770] = 13;
// bram[45771] = 5;
// bram[45772] = 1;
// bram[45773] = 0;
// bram[45774] = 3;
// bram[45775] = 9;
// bram[45776] = 19;
// bram[45777] = 33;
// bram[45778] = 49;
// bram[45779] = 67;
// bram[45780] = 87;
// bram[45781] = 109;
// bram[45782] = 130;
// bram[45783] = 152;
// bram[45784] = 173;
// bram[45785] = 193;
// bram[45786] = 210;
// bram[45787] = 226;
// bram[45788] = 238;
// bram[45789] = 247;
// bram[45790] = 252;
// bram[45791] = 253;
// bram[45792] = 251;
// bram[45793] = 245;
// bram[45794] = 236;
// bram[45795] = 223;
// bram[45796] = 207;
// bram[45797] = 189;
// bram[45798] = 170;
// bram[45799] = 148;
// bram[45800] = 127;
// bram[45801] = 105;
// bram[45802] = 83;
// bram[45803] = 64;
// bram[45804] = 46;
// bram[45805] = 30;
// bram[45806] = 17;
// bram[45807] = 8;
// bram[45808] = 2;
// bram[45809] = 0;
// bram[45810] = 1;
// bram[45811] = 6;
// bram[45812] = 15;
// bram[45813] = 27;
// bram[45814] = 43;
// bram[45815] = 60;
// bram[45816] = 80;
// bram[45817] = 101;
// bram[45818] = 123;
// bram[45819] = 144;
// bram[45820] = 166;
// bram[45821] = 186;
// bram[45822] = 204;
// bram[45823] = 220;
// bram[45824] = 234;
// bram[45825] = 244;
// bram[45826] = 250;
// bram[45827] = 253;
// bram[45828] = 252;
// bram[45829] = 248;
// bram[45830] = 240;
// bram[45831] = 228;
// bram[45832] = 213;
// bram[45833] = 196;
// bram[45834] = 177;
// bram[45835] = 156;
// bram[45836] = 134;
// bram[45837] = 113;
// bram[45838] = 91;
// bram[45839] = 71;
// bram[45840] = 52;
// bram[45841] = 35;
// bram[45842] = 21;
// bram[45843] = 11;
// bram[45844] = 3;
// bram[45845] = 0;
// bram[45846] = 0;
// bram[45847] = 4;
// bram[45848] = 12;
// bram[45849] = 23;
// bram[45850] = 37;
// bram[45851] = 53;
// bram[45852] = 72;
// bram[45853] = 93;
// bram[45854] = 115;
// bram[45855] = 136;
// bram[45856] = 158;
// bram[45857] = 179;
// bram[45858] = 198;
// bram[45859] = 215;
// bram[45860] = 229;
// bram[45861] = 241;
// bram[45862] = 248;
// bram[45863] = 253;
// bram[45864] = 253;
// bram[45865] = 250;
// bram[45866] = 243;
// bram[45867] = 233;
// bram[45868] = 219;
// bram[45869] = 203;
// bram[45870] = 184;
// bram[45871] = 164;
// bram[45872] = 142;
// bram[45873] = 121;
// bram[45874] = 99;
// bram[45875] = 78;
// bram[45876] = 58;
// bram[45877] = 41;
// bram[45878] = 26;
// bram[45879] = 14;
// bram[45880] = 6;
// bram[45881] = 1;
// bram[45882] = 0;
// bram[45883] = 2;
// bram[45884] = 8;
// bram[45885] = 18;
// bram[45886] = 31;
// bram[45887] = 47;
// bram[45888] = 65;
// bram[45889] = 85;
// bram[45890] = 107;
// bram[45891] = 128;
// bram[45892] = 150;
// bram[45893] = 171;
// bram[45894] = 191;
// bram[45895] = 209;
// bram[45896] = 224;
// bram[45897] = 237;
// bram[45898] = 246;
// bram[45899] = 252;
// bram[45900] = 254;
// bram[45901] = 252;
// bram[45902] = 246;
// bram[45903] = 237;
// bram[45904] = 224;
// bram[45905] = 209;
// bram[45906] = 191;
// bram[45907] = 171;
// bram[45908] = 150;
// bram[45909] = 128;
// bram[45910] = 107;
// bram[45911] = 85;
// bram[45912] = 65;
// bram[45913] = 47;
// bram[45914] = 31;
// bram[45915] = 18;
// bram[45916] = 8;
// bram[45917] = 2;
// bram[45918] = 0;
// bram[45919] = 1;
// bram[45920] = 6;
// bram[45921] = 14;
// bram[45922] = 26;
// bram[45923] = 41;
// bram[45924] = 58;
// bram[45925] = 78;
// bram[45926] = 99;
// bram[45927] = 121;
// bram[45928] = 142;
// bram[45929] = 164;
// bram[45930] = 184;
// bram[45931] = 203;
// bram[45932] = 219;
// bram[45933] = 233;
// bram[45934] = 243;
// bram[45935] = 250;
// bram[45936] = 253;
// bram[45937] = 253;
// bram[45938] = 248;
// bram[45939] = 241;
// bram[45940] = 229;
// bram[45941] = 215;
// bram[45942] = 198;
// bram[45943] = 179;
// bram[45944] = 158;
// bram[45945] = 136;
// bram[45946] = 115;
// bram[45947] = 93;
// bram[45948] = 72;
// bram[45949] = 53;
// bram[45950] = 37;
// bram[45951] = 23;
// bram[45952] = 12;
// bram[45953] = 4;
// bram[45954] = 0;
// bram[45955] = 0;
// bram[45956] = 3;
// bram[45957] = 11;
// bram[45958] = 21;
// bram[45959] = 35;
// bram[45960] = 52;
// bram[45961] = 71;
// bram[45962] = 91;
// bram[45963] = 113;
// bram[45964] = 134;
// bram[45965] = 156;
// bram[45966] = 177;
// bram[45967] = 196;
// bram[45968] = 213;
// bram[45969] = 228;
// bram[45970] = 240;
// bram[45971] = 248;
// bram[45972] = 252;
// bram[45973] = 253;
// bram[45974] = 250;
// bram[45975] = 244;
// bram[45976] = 234;
// bram[45977] = 220;
// bram[45978] = 204;
// bram[45979] = 186;
// bram[45980] = 166;
// bram[45981] = 144;
// bram[45982] = 123;
// bram[45983] = 101;
// bram[45984] = 80;
// bram[45985] = 60;
// bram[45986] = 43;
// bram[45987] = 27;
// bram[45988] = 15;
// bram[45989] = 6;
// bram[45990] = 1;
// bram[45991] = 0;
// bram[45992] = 2;
// bram[45993] = 8;
// bram[45994] = 17;
// bram[45995] = 30;
// bram[45996] = 46;
// bram[45997] = 64;
// bram[45998] = 83;
// bram[45999] = 105;
// bram[46000] = 127;
// bram[46001] = 148;
// bram[46002] = 170;
// bram[46003] = 189;
// bram[46004] = 207;
// bram[46005] = 223;
// bram[46006] = 236;
// bram[46007] = 245;
// bram[46008] = 251;
// bram[46009] = 253;
// bram[46010] = 252;
// bram[46011] = 247;
// bram[46012] = 238;
// bram[46013] = 226;
// bram[46014] = 210;
// bram[46015] = 193;
// bram[46016] = 173;
// bram[46017] = 152;
// bram[46018] = 130;
// bram[46019] = 109;
// bram[46020] = 87;
// bram[46021] = 67;
// bram[46022] = 49;
// bram[46023] = 33;
// bram[46024] = 19;
// bram[46025] = 9;
// bram[46026] = 3;
// bram[46027] = 0;
// bram[46028] = 1;
// bram[46029] = 5;
// bram[46030] = 13;
// bram[46031] = 25;
// bram[46032] = 40;
// bram[46033] = 57;
// bram[46034] = 76;
// bram[46035] = 97;
// bram[46036] = 119;
// bram[46037] = 140;
// bram[46038] = 162;
// bram[46039] = 182;
// bram[46040] = 201;
// bram[46041] = 218;
// bram[46042] = 232;
// bram[46043] = 242;
// bram[46044] = 250;
// bram[46045] = 253;
// bram[46046] = 253;
// bram[46047] = 249;
// bram[46048] = 241;
// bram[46049] = 230;
// bram[46050] = 216;
// bram[46051] = 200;
// bram[46052] = 181;
// bram[46053] = 160;
// bram[46054] = 138;
// bram[46055] = 117;
// bram[46056] = 95;
// bram[46057] = 74;
// bram[46058] = 55;
// bram[46059] = 38;
// bram[46060] = 24;
// bram[46061] = 12;
// bram[46062] = 5;
// bram[46063] = 0;
// bram[46064] = 0;
// bram[46065] = 3;
// bram[46066] = 10;
// bram[46067] = 20;
// bram[46068] = 34;
// bram[46069] = 50;
// bram[46070] = 69;
// bram[46071] = 89;
// bram[46072] = 111;
// bram[46073] = 132;
// bram[46074] = 154;
// bram[46075] = 175;
// bram[46076] = 195;
// bram[46077] = 212;
// bram[46078] = 227;
// bram[46079] = 239;
// bram[46080] = 247;
// bram[46081] = 252;
// bram[46082] = 253;
// bram[46083] = 251;
// bram[46084] = 245;
// bram[46085] = 235;
// bram[46086] = 222;
// bram[46087] = 206;
// bram[46088] = 188;
// bram[46089] = 168;
// bram[46090] = 146;
// bram[46091] = 125;
// bram[46092] = 103;
// bram[46093] = 82;
// bram[46094] = 62;
// bram[46095] = 44;
// bram[46096] = 29;
// bram[46097] = 16;
// bram[46098] = 7;
// bram[46099] = 1;
// bram[46100] = 0;
// bram[46101] = 1;
// bram[46102] = 7;
// bram[46103] = 16;
// bram[46104] = 29;
// bram[46105] = 44;
// bram[46106] = 62;
// bram[46107] = 82;
// bram[46108] = 103;
// bram[46109] = 125;
// bram[46110] = 146;
// bram[46111] = 168;
// bram[46112] = 188;
// bram[46113] = 206;
// bram[46114] = 222;
// bram[46115] = 235;
// bram[46116] = 245;
// bram[46117] = 251;
// bram[46118] = 253;
// bram[46119] = 252;
// bram[46120] = 247;
// bram[46121] = 239;
// bram[46122] = 227;
// bram[46123] = 212;
// bram[46124] = 195;
// bram[46125] = 175;
// bram[46126] = 154;
// bram[46127] = 132;
// bram[46128] = 111;
// bram[46129] = 89;
// bram[46130] = 69;
// bram[46131] = 50;
// bram[46132] = 34;
// bram[46133] = 20;
// bram[46134] = 10;
// bram[46135] = 3;
// bram[46136] = 0;
// bram[46137] = 0;
// bram[46138] = 5;
// bram[46139] = 12;
// bram[46140] = 24;
// bram[46141] = 38;
// bram[46142] = 55;
// bram[46143] = 74;
// bram[46144] = 95;
// bram[46145] = 117;
// bram[46146] = 138;
// bram[46147] = 160;
// bram[46148] = 181;
// bram[46149] = 200;
// bram[46150] = 216;
// bram[46151] = 230;
// bram[46152] = 241;
// bram[46153] = 249;
// bram[46154] = 253;
// bram[46155] = 253;
// bram[46156] = 250;
// bram[46157] = 242;
// bram[46158] = 232;
// bram[46159] = 218;
// bram[46160] = 201;
// bram[46161] = 182;
// bram[46162] = 162;
// bram[46163] = 140;
// bram[46164] = 119;
// bram[46165] = 97;
// bram[46166] = 76;
// bram[46167] = 57;
// bram[46168] = 40;
// bram[46169] = 25;
// bram[46170] = 13;
// bram[46171] = 5;
// bram[46172] = 1;
// bram[46173] = 0;
// bram[46174] = 3;
// bram[46175] = 9;
// bram[46176] = 19;
// bram[46177] = 33;
// bram[46178] = 49;
// bram[46179] = 67;
// bram[46180] = 87;
// bram[46181] = 109;
// bram[46182] = 130;
// bram[46183] = 152;
// bram[46184] = 173;
// bram[46185] = 193;
// bram[46186] = 210;
// bram[46187] = 226;
// bram[46188] = 238;
// bram[46189] = 247;
// bram[46190] = 252;
// bram[46191] = 253;
// bram[46192] = 251;
// bram[46193] = 245;
// bram[46194] = 236;
// bram[46195] = 223;
// bram[46196] = 207;
// bram[46197] = 189;
// bram[46198] = 170;
// bram[46199] = 148;
// bram[46200] = 126;
// bram[46201] = 105;
// bram[46202] = 83;
// bram[46203] = 64;
// bram[46204] = 46;
// bram[46205] = 30;
// bram[46206] = 17;
// bram[46207] = 8;
// bram[46208] = 2;
// bram[46209] = 0;
// bram[46210] = 1;
// bram[46211] = 6;
// bram[46212] = 15;
// bram[46213] = 27;
// bram[46214] = 43;
// bram[46215] = 60;
// bram[46216] = 80;
// bram[46217] = 101;
// bram[46218] = 123;
// bram[46219] = 144;
// bram[46220] = 166;
// bram[46221] = 186;
// bram[46222] = 204;
// bram[46223] = 220;
// bram[46224] = 234;
// bram[46225] = 244;
// bram[46226] = 250;
// bram[46227] = 253;
// bram[46228] = 252;
// bram[46229] = 248;
// bram[46230] = 240;
// bram[46231] = 228;
// bram[46232] = 213;
// bram[46233] = 196;
// bram[46234] = 177;
// bram[46235] = 156;
// bram[46236] = 134;
// bram[46237] = 113;
// bram[46238] = 91;
// bram[46239] = 71;
// bram[46240] = 52;
// bram[46241] = 35;
// bram[46242] = 21;
// bram[46243] = 11;
// bram[46244] = 3;
// bram[46245] = 0;
// bram[46246] = 0;
// bram[46247] = 4;
// bram[46248] = 12;
// bram[46249] = 23;
// bram[46250] = 37;
// bram[46251] = 53;
// bram[46252] = 72;
// bram[46253] = 93;
// bram[46254] = 115;
// bram[46255] = 136;
// bram[46256] = 158;
// bram[46257] = 179;
// bram[46258] = 198;
// bram[46259] = 215;
// bram[46260] = 229;
// bram[46261] = 241;
// bram[46262] = 248;
// bram[46263] = 253;
// bram[46264] = 253;
// bram[46265] = 250;
// bram[46266] = 243;
// bram[46267] = 233;
// bram[46268] = 219;
// bram[46269] = 203;
// bram[46270] = 184;
// bram[46271] = 164;
// bram[46272] = 142;
// bram[46273] = 121;
// bram[46274] = 99;
// bram[46275] = 78;
// bram[46276] = 58;
// bram[46277] = 41;
// bram[46278] = 26;
// bram[46279] = 14;
// bram[46280] = 6;
// bram[46281] = 1;
// bram[46282] = 0;
// bram[46283] = 2;
// bram[46284] = 8;
// bram[46285] = 18;
// bram[46286] = 31;
// bram[46287] = 47;
// bram[46288] = 65;
// bram[46289] = 85;
// bram[46290] = 107;
// bram[46291] = 128;
// bram[46292] = 150;
// bram[46293] = 171;
// bram[46294] = 191;
// bram[46295] = 209;
// bram[46296] = 224;
// bram[46297] = 237;
// bram[46298] = 246;
// bram[46299] = 252;
// bram[46300] = 254;
// bram[46301] = 252;
// bram[46302] = 246;
// bram[46303] = 237;
// bram[46304] = 224;
// bram[46305] = 209;
// bram[46306] = 191;
// bram[46307] = 171;
// bram[46308] = 150;
// bram[46309] = 128;
// bram[46310] = 107;
// bram[46311] = 85;
// bram[46312] = 65;
// bram[46313] = 47;
// bram[46314] = 31;
// bram[46315] = 18;
// bram[46316] = 8;
// bram[46317] = 2;
// bram[46318] = 0;
// bram[46319] = 1;
// bram[46320] = 6;
// bram[46321] = 14;
// bram[46322] = 26;
// bram[46323] = 41;
// bram[46324] = 58;
// bram[46325] = 78;
// bram[46326] = 99;
// bram[46327] = 121;
// bram[46328] = 142;
// bram[46329] = 164;
// bram[46330] = 184;
// bram[46331] = 203;
// bram[46332] = 219;
// bram[46333] = 233;
// bram[46334] = 243;
// bram[46335] = 250;
// bram[46336] = 253;
// bram[46337] = 253;
// bram[46338] = 248;
// bram[46339] = 241;
// bram[46340] = 229;
// bram[46341] = 215;
// bram[46342] = 198;
// bram[46343] = 179;
// bram[46344] = 158;
// bram[46345] = 136;
// bram[46346] = 115;
// bram[46347] = 93;
// bram[46348] = 72;
// bram[46349] = 53;
// bram[46350] = 37;
// bram[46351] = 23;
// bram[46352] = 12;
// bram[46353] = 4;
// bram[46354] = 0;
// bram[46355] = 0;
// bram[46356] = 3;
// bram[46357] = 11;
// bram[46358] = 21;
// bram[46359] = 35;
// bram[46360] = 52;
// bram[46361] = 71;
// bram[46362] = 91;
// bram[46363] = 113;
// bram[46364] = 134;
// bram[46365] = 156;
// bram[46366] = 177;
// bram[46367] = 196;
// bram[46368] = 213;
// bram[46369] = 228;
// bram[46370] = 240;
// bram[46371] = 248;
// bram[46372] = 252;
// bram[46373] = 253;
// bram[46374] = 250;
// bram[46375] = 244;
// bram[46376] = 234;
// bram[46377] = 220;
// bram[46378] = 204;
// bram[46379] = 186;
// bram[46380] = 166;
// bram[46381] = 144;
// bram[46382] = 123;
// bram[46383] = 101;
// bram[46384] = 80;
// bram[46385] = 60;
// bram[46386] = 43;
// bram[46387] = 27;
// bram[46388] = 15;
// bram[46389] = 6;
// bram[46390] = 1;
// bram[46391] = 0;
// bram[46392] = 2;
// bram[46393] = 8;
// bram[46394] = 17;
// bram[46395] = 30;
// bram[46396] = 46;
// bram[46397] = 64;
// bram[46398] = 83;
// bram[46399] = 105;
// bram[46400] = 127;
// bram[46401] = 148;
// bram[46402] = 170;
// bram[46403] = 189;
// bram[46404] = 207;
// bram[46405] = 223;
// bram[46406] = 236;
// bram[46407] = 245;
// bram[46408] = 251;
// bram[46409] = 253;
// bram[46410] = 252;
// bram[46411] = 247;
// bram[46412] = 238;
// bram[46413] = 226;
// bram[46414] = 210;
// bram[46415] = 193;
// bram[46416] = 173;
// bram[46417] = 152;
// bram[46418] = 130;
// bram[46419] = 109;
// bram[46420] = 87;
// bram[46421] = 67;
// bram[46422] = 49;
// bram[46423] = 33;
// bram[46424] = 19;
// bram[46425] = 9;
// bram[46426] = 3;
// bram[46427] = 0;
// bram[46428] = 1;
// bram[46429] = 5;
// bram[46430] = 13;
// bram[46431] = 25;
// bram[46432] = 40;
// bram[46433] = 57;
// bram[46434] = 76;
// bram[46435] = 97;
// bram[46436] = 119;
// bram[46437] = 140;
// bram[46438] = 162;
// bram[46439] = 182;
// bram[46440] = 201;
// bram[46441] = 218;
// bram[46442] = 232;
// bram[46443] = 242;
// bram[46444] = 250;
// bram[46445] = 253;
// bram[46446] = 253;
// bram[46447] = 249;
// bram[46448] = 241;
// bram[46449] = 230;
// bram[46450] = 216;
// bram[46451] = 200;
// bram[46452] = 181;
// bram[46453] = 160;
// bram[46454] = 138;
// bram[46455] = 117;
// bram[46456] = 95;
// bram[46457] = 74;
// bram[46458] = 55;
// bram[46459] = 38;
// bram[46460] = 24;
// bram[46461] = 12;
// bram[46462] = 5;
// bram[46463] = 0;
// bram[46464] = 0;
// bram[46465] = 3;
// bram[46466] = 10;
// bram[46467] = 20;
// bram[46468] = 34;
// bram[46469] = 50;
// bram[46470] = 69;
// bram[46471] = 89;
// bram[46472] = 111;
// bram[46473] = 132;
// bram[46474] = 154;
// bram[46475] = 175;
// bram[46476] = 195;
// bram[46477] = 212;
// bram[46478] = 227;
// bram[46479] = 239;
// bram[46480] = 247;
// bram[46481] = 252;
// bram[46482] = 253;
// bram[46483] = 251;
// bram[46484] = 245;
// bram[46485] = 235;
// bram[46486] = 222;
// bram[46487] = 206;
// bram[46488] = 188;
// bram[46489] = 168;
// bram[46490] = 146;
// bram[46491] = 125;
// bram[46492] = 103;
// bram[46493] = 82;
// bram[46494] = 62;
// bram[46495] = 44;
// bram[46496] = 29;
// bram[46497] = 16;
// bram[46498] = 7;
// bram[46499] = 1;
// bram[46500] = 0;
// bram[46501] = 1;
// bram[46502] = 7;
// bram[46503] = 16;
// bram[46504] = 29;
// bram[46505] = 44;
// bram[46506] = 62;
// bram[46507] = 82;
// bram[46508] = 103;
// bram[46509] = 125;
// bram[46510] = 146;
// bram[46511] = 168;
// bram[46512] = 188;
// bram[46513] = 206;
// bram[46514] = 222;
// bram[46515] = 235;
// bram[46516] = 245;
// bram[46517] = 251;
// bram[46518] = 253;
// bram[46519] = 252;
// bram[46520] = 247;
// bram[46521] = 239;
// bram[46522] = 227;
// bram[46523] = 212;
// bram[46524] = 195;
// bram[46525] = 175;
// bram[46526] = 154;
// bram[46527] = 132;
// bram[46528] = 111;
// bram[46529] = 89;
// bram[46530] = 69;
// bram[46531] = 50;
// bram[46532] = 34;
// bram[46533] = 20;
// bram[46534] = 10;
// bram[46535] = 3;
// bram[46536] = 0;
// bram[46537] = 0;
// bram[46538] = 5;
// bram[46539] = 12;
// bram[46540] = 24;
// bram[46541] = 38;
// bram[46542] = 55;
// bram[46543] = 74;
// bram[46544] = 95;
// bram[46545] = 117;
// bram[46546] = 138;
// bram[46547] = 160;
// bram[46548] = 181;
// bram[46549] = 200;
// bram[46550] = 216;
// bram[46551] = 230;
// bram[46552] = 241;
// bram[46553] = 249;
// bram[46554] = 253;
// bram[46555] = 253;
// bram[46556] = 250;
// bram[46557] = 242;
// bram[46558] = 232;
// bram[46559] = 218;
// bram[46560] = 201;
// bram[46561] = 182;
// bram[46562] = 162;
// bram[46563] = 140;
// bram[46564] = 119;
// bram[46565] = 97;
// bram[46566] = 76;
// bram[46567] = 57;
// bram[46568] = 40;
// bram[46569] = 25;
// bram[46570] = 13;
// bram[46571] = 5;
// bram[46572] = 1;
// bram[46573] = 0;
// bram[46574] = 3;
// bram[46575] = 9;
// bram[46576] = 19;
// bram[46577] = 33;
// bram[46578] = 49;
// bram[46579] = 67;
// bram[46580] = 87;
// bram[46581] = 109;
// bram[46582] = 130;
// bram[46583] = 152;
// bram[46584] = 173;
// bram[46585] = 193;
// bram[46586] = 210;
// bram[46587] = 226;
// bram[46588] = 238;
// bram[46589] = 247;
// bram[46590] = 252;
// bram[46591] = 253;
// bram[46592] = 251;
// bram[46593] = 245;
// bram[46594] = 236;
// bram[46595] = 223;
// bram[46596] = 207;
// bram[46597] = 189;
// bram[46598] = 170;
// bram[46599] = 148;
// bram[46600] = 126;
// bram[46601] = 105;
// bram[46602] = 83;
// bram[46603] = 64;
// bram[46604] = 46;
// bram[46605] = 30;
// bram[46606] = 17;
// bram[46607] = 8;
// bram[46608] = 2;
// bram[46609] = 0;
// bram[46610] = 1;
// bram[46611] = 6;
// bram[46612] = 15;
// bram[46613] = 27;
// bram[46614] = 43;
// bram[46615] = 60;
// bram[46616] = 80;
// bram[46617] = 101;
// bram[46618] = 123;
// bram[46619] = 144;
// bram[46620] = 166;
// bram[46621] = 186;
// bram[46622] = 204;
// bram[46623] = 220;
// bram[46624] = 234;
// bram[46625] = 244;
// bram[46626] = 250;
// bram[46627] = 253;
// bram[46628] = 252;
// bram[46629] = 248;
// bram[46630] = 240;
// bram[46631] = 228;
// bram[46632] = 213;
// bram[46633] = 196;
// bram[46634] = 177;
// bram[46635] = 156;
// bram[46636] = 134;
// bram[46637] = 113;
// bram[46638] = 91;
// bram[46639] = 71;
// bram[46640] = 52;
// bram[46641] = 35;
// bram[46642] = 21;
// bram[46643] = 11;
// bram[46644] = 3;
// bram[46645] = 0;
// bram[46646] = 0;
// bram[46647] = 4;
// bram[46648] = 12;
// bram[46649] = 23;
// bram[46650] = 37;
// bram[46651] = 53;
// bram[46652] = 72;
// bram[46653] = 93;
// bram[46654] = 115;
// bram[46655] = 136;
// bram[46656] = 158;
// bram[46657] = 179;
// bram[46658] = 198;
// bram[46659] = 215;
// bram[46660] = 229;
// bram[46661] = 241;
// bram[46662] = 248;
// bram[46663] = 253;
// bram[46664] = 253;
// bram[46665] = 250;
// bram[46666] = 243;
// bram[46667] = 233;
// bram[46668] = 219;
// bram[46669] = 203;
// bram[46670] = 184;
// bram[46671] = 164;
// bram[46672] = 142;
// bram[46673] = 121;
// bram[46674] = 99;
// bram[46675] = 78;
// bram[46676] = 58;
// bram[46677] = 41;
// bram[46678] = 26;
// bram[46679] = 14;
// bram[46680] = 6;
// bram[46681] = 1;
// bram[46682] = 0;
// bram[46683] = 2;
// bram[46684] = 8;
// bram[46685] = 18;
// bram[46686] = 31;
// bram[46687] = 47;
// bram[46688] = 65;
// bram[46689] = 85;
// bram[46690] = 107;
// bram[46691] = 128;
// bram[46692] = 150;
// bram[46693] = 171;
// bram[46694] = 191;
// bram[46695] = 209;
// bram[46696] = 224;
// bram[46697] = 237;
// bram[46698] = 246;
// bram[46699] = 252;
// bram[46700] = 254;
// bram[46701] = 252;
// bram[46702] = 246;
// bram[46703] = 237;
// bram[46704] = 224;
// bram[46705] = 209;
// bram[46706] = 191;
// bram[46707] = 171;
// bram[46708] = 150;
// bram[46709] = 128;
// bram[46710] = 107;
// bram[46711] = 85;
// bram[46712] = 65;
// bram[46713] = 47;
// bram[46714] = 31;
// bram[46715] = 18;
// bram[46716] = 8;
// bram[46717] = 2;
// bram[46718] = 0;
// bram[46719] = 1;
// bram[46720] = 6;
// bram[46721] = 14;
// bram[46722] = 26;
// bram[46723] = 41;
// bram[46724] = 58;
// bram[46725] = 78;
// bram[46726] = 99;
// bram[46727] = 121;
// bram[46728] = 142;
// bram[46729] = 164;
// bram[46730] = 184;
// bram[46731] = 203;
// bram[46732] = 219;
// bram[46733] = 233;
// bram[46734] = 243;
// bram[46735] = 250;
// bram[46736] = 253;
// bram[46737] = 253;
// bram[46738] = 248;
// bram[46739] = 241;
// bram[46740] = 229;
// bram[46741] = 215;
// bram[46742] = 198;
// bram[46743] = 179;
// bram[46744] = 158;
// bram[46745] = 136;
// bram[46746] = 115;
// bram[46747] = 93;
// bram[46748] = 72;
// bram[46749] = 53;
// bram[46750] = 37;
// bram[46751] = 23;
// bram[46752] = 12;
// bram[46753] = 4;
// bram[46754] = 0;
// bram[46755] = 0;
// bram[46756] = 3;
// bram[46757] = 11;
// bram[46758] = 21;
// bram[46759] = 35;
// bram[46760] = 52;
// bram[46761] = 71;
// bram[46762] = 91;
// bram[46763] = 113;
// bram[46764] = 134;
// bram[46765] = 156;
// bram[46766] = 177;
// bram[46767] = 196;
// bram[46768] = 213;
// bram[46769] = 228;
// bram[46770] = 240;
// bram[46771] = 248;
// bram[46772] = 252;
// bram[46773] = 253;
// bram[46774] = 250;
// bram[46775] = 244;
// bram[46776] = 234;
// bram[46777] = 220;
// bram[46778] = 204;
// bram[46779] = 186;
// bram[46780] = 166;
// bram[46781] = 144;
// bram[46782] = 123;
// bram[46783] = 101;
// bram[46784] = 80;
// bram[46785] = 60;
// bram[46786] = 43;
// bram[46787] = 27;
// bram[46788] = 15;
// bram[46789] = 6;
// bram[46790] = 1;
// bram[46791] = 0;
// bram[46792] = 2;
// bram[46793] = 8;
// bram[46794] = 17;
// bram[46795] = 30;
// bram[46796] = 46;
// bram[46797] = 64;
// bram[46798] = 83;
// bram[46799] = 105;
// bram[46800] = 127;
// bram[46801] = 148;
// bram[46802] = 170;
// bram[46803] = 189;
// bram[46804] = 207;
// bram[46805] = 223;
// bram[46806] = 236;
// bram[46807] = 245;
// bram[46808] = 251;
// bram[46809] = 253;
// bram[46810] = 252;
// bram[46811] = 247;
// bram[46812] = 238;
// bram[46813] = 226;
// bram[46814] = 210;
// bram[46815] = 193;
// bram[46816] = 173;
// bram[46817] = 152;
// bram[46818] = 130;
// bram[46819] = 109;
// bram[46820] = 87;
// bram[46821] = 67;
// bram[46822] = 49;
// bram[46823] = 33;
// bram[46824] = 19;
// bram[46825] = 9;
// bram[46826] = 3;
// bram[46827] = 0;
// bram[46828] = 1;
// bram[46829] = 5;
// bram[46830] = 13;
// bram[46831] = 25;
// bram[46832] = 40;
// bram[46833] = 57;
// bram[46834] = 76;
// bram[46835] = 97;
// bram[46836] = 119;
// bram[46837] = 140;
// bram[46838] = 162;
// bram[46839] = 182;
// bram[46840] = 201;
// bram[46841] = 218;
// bram[46842] = 232;
// bram[46843] = 242;
// bram[46844] = 250;
// bram[46845] = 253;
// bram[46846] = 253;
// bram[46847] = 249;
// bram[46848] = 241;
// bram[46849] = 230;
// bram[46850] = 216;
// bram[46851] = 200;
// bram[46852] = 181;
// bram[46853] = 160;
// bram[46854] = 138;
// bram[46855] = 117;
// bram[46856] = 95;
// bram[46857] = 74;
// bram[46858] = 55;
// bram[46859] = 38;
// bram[46860] = 24;
// bram[46861] = 12;
// bram[46862] = 5;
// bram[46863] = 0;
// bram[46864] = 0;
// bram[46865] = 3;
// bram[46866] = 10;
// bram[46867] = 20;
// bram[46868] = 34;
// bram[46869] = 50;
// bram[46870] = 69;
// bram[46871] = 89;
// bram[46872] = 111;
// bram[46873] = 132;
// bram[46874] = 154;
// bram[46875] = 175;
// bram[46876] = 195;
// bram[46877] = 212;
// bram[46878] = 227;
// bram[46879] = 239;
// bram[46880] = 247;
// bram[46881] = 252;
// bram[46882] = 253;
// bram[46883] = 251;
// bram[46884] = 245;
// bram[46885] = 235;
// bram[46886] = 222;
// bram[46887] = 206;
// bram[46888] = 188;
// bram[46889] = 168;
// bram[46890] = 146;
// bram[46891] = 125;
// bram[46892] = 103;
// bram[46893] = 82;
// bram[46894] = 62;
// bram[46895] = 44;
// bram[46896] = 29;
// bram[46897] = 16;
// bram[46898] = 7;
// bram[46899] = 1;
// bram[46900] = 0;
// bram[46901] = 1;
// bram[46902] = 7;
// bram[46903] = 16;
// bram[46904] = 29;
// bram[46905] = 44;
// bram[46906] = 62;
// bram[46907] = 82;
// bram[46908] = 103;
// bram[46909] = 125;
// bram[46910] = 146;
// bram[46911] = 168;
// bram[46912] = 188;
// bram[46913] = 206;
// bram[46914] = 222;
// bram[46915] = 235;
// bram[46916] = 245;
// bram[46917] = 251;
// bram[46918] = 253;
// bram[46919] = 252;
// bram[46920] = 247;
// bram[46921] = 239;
// bram[46922] = 227;
// bram[46923] = 212;
// bram[46924] = 195;
// bram[46925] = 175;
// bram[46926] = 154;
// bram[46927] = 132;
// bram[46928] = 111;
// bram[46929] = 89;
// bram[46930] = 69;
// bram[46931] = 50;
// bram[46932] = 34;
// bram[46933] = 20;
// bram[46934] = 10;
// bram[46935] = 3;
// bram[46936] = 0;
// bram[46937] = 0;
// bram[46938] = 5;
// bram[46939] = 12;
// bram[46940] = 24;
// bram[46941] = 38;
// bram[46942] = 55;
// bram[46943] = 74;
// bram[46944] = 95;
// bram[46945] = 117;
// bram[46946] = 138;
// bram[46947] = 160;
// bram[46948] = 181;
// bram[46949] = 200;
// bram[46950] = 216;
// bram[46951] = 230;
// bram[46952] = 241;
// bram[46953] = 249;
// bram[46954] = 253;
// bram[46955] = 253;
// bram[46956] = 250;
// bram[46957] = 242;
// bram[46958] = 232;
// bram[46959] = 218;
// bram[46960] = 201;
// bram[46961] = 182;
// bram[46962] = 162;
// bram[46963] = 140;
// bram[46964] = 119;
// bram[46965] = 97;
// bram[46966] = 76;
// bram[46967] = 57;
// bram[46968] = 40;
// bram[46969] = 25;
// bram[46970] = 13;
// bram[46971] = 5;
// bram[46972] = 1;
// bram[46973] = 0;
// bram[46974] = 3;
// bram[46975] = 9;
// bram[46976] = 19;
// bram[46977] = 33;
// bram[46978] = 49;
// bram[46979] = 67;
// bram[46980] = 87;
// bram[46981] = 109;
// bram[46982] = 130;
// bram[46983] = 152;
// bram[46984] = 173;
// bram[46985] = 193;
// bram[46986] = 210;
// bram[46987] = 226;
// bram[46988] = 238;
// bram[46989] = 247;
// bram[46990] = 252;
// bram[46991] = 253;
// bram[46992] = 251;
// bram[46993] = 245;
// bram[46994] = 236;
// bram[46995] = 223;
// bram[46996] = 207;
// bram[46997] = 189;
// bram[46998] = 170;
// bram[46999] = 148;
// bram[47000] = 126;
// bram[47001] = 105;
// bram[47002] = 83;
// bram[47003] = 64;
// bram[47004] = 46;
// bram[47005] = 30;
// bram[47006] = 17;
// bram[47007] = 8;
// bram[47008] = 2;
// bram[47009] = 0;
// bram[47010] = 1;
// bram[47011] = 6;
// bram[47012] = 15;
// bram[47013] = 27;
// bram[47014] = 43;
// bram[47015] = 60;
// bram[47016] = 80;
// bram[47017] = 101;
// bram[47018] = 123;
// bram[47019] = 144;
// bram[47020] = 166;
// bram[47021] = 186;
// bram[47022] = 204;
// bram[47023] = 220;
// bram[47024] = 234;
// bram[47025] = 244;
// bram[47026] = 250;
// bram[47027] = 253;
// bram[47028] = 252;
// bram[47029] = 248;
// bram[47030] = 240;
// bram[47031] = 228;
// bram[47032] = 213;
// bram[47033] = 196;
// bram[47034] = 177;
// bram[47035] = 156;
// bram[47036] = 134;
// bram[47037] = 113;
// bram[47038] = 91;
// bram[47039] = 71;
// bram[47040] = 52;
// bram[47041] = 35;
// bram[47042] = 21;
// bram[47043] = 11;
// bram[47044] = 3;
// bram[47045] = 0;
// bram[47046] = 0;
// bram[47047] = 4;
// bram[47048] = 12;
// bram[47049] = 23;
// bram[47050] = 37;
// bram[47051] = 53;
// bram[47052] = 72;
// bram[47053] = 93;
// bram[47054] = 115;
// bram[47055] = 136;
// bram[47056] = 158;
// bram[47057] = 179;
// bram[47058] = 198;
// bram[47059] = 215;
// bram[47060] = 229;
// bram[47061] = 241;
// bram[47062] = 248;
// bram[47063] = 253;
// bram[47064] = 253;
// bram[47065] = 250;
// bram[47066] = 243;
// bram[47067] = 233;
// bram[47068] = 219;
// bram[47069] = 203;
// bram[47070] = 184;
// bram[47071] = 164;
// bram[47072] = 142;
// bram[47073] = 121;
// bram[47074] = 99;
// bram[47075] = 78;
// bram[47076] = 58;
// bram[47077] = 41;
// bram[47078] = 26;
// bram[47079] = 14;
// bram[47080] = 6;
// bram[47081] = 1;
// bram[47082] = 0;
// bram[47083] = 2;
// bram[47084] = 8;
// bram[47085] = 18;
// bram[47086] = 31;
// bram[47087] = 47;
// bram[47088] = 65;
// bram[47089] = 85;
// bram[47090] = 107;
// bram[47091] = 128;
// bram[47092] = 150;
// bram[47093] = 171;
// bram[47094] = 191;
// bram[47095] = 209;
// bram[47096] = 224;
// bram[47097] = 237;
// bram[47098] = 246;
// bram[47099] = 252;
// bram[47100] = 254;
// bram[47101] = 252;
// bram[47102] = 246;
// bram[47103] = 237;
// bram[47104] = 224;
// bram[47105] = 209;
// bram[47106] = 191;
// bram[47107] = 171;
// bram[47108] = 150;
// bram[47109] = 128;
// bram[47110] = 107;
// bram[47111] = 85;
// bram[47112] = 65;
// bram[47113] = 47;
// bram[47114] = 31;
// bram[47115] = 18;
// bram[47116] = 8;
// bram[47117] = 2;
// bram[47118] = 0;
// bram[47119] = 1;
// bram[47120] = 6;
// bram[47121] = 14;
// bram[47122] = 26;
// bram[47123] = 41;
// bram[47124] = 58;
// bram[47125] = 78;
// bram[47126] = 99;
// bram[47127] = 121;
// bram[47128] = 142;
// bram[47129] = 164;
// bram[47130] = 184;
// bram[47131] = 203;
// bram[47132] = 219;
// bram[47133] = 233;
// bram[47134] = 243;
// bram[47135] = 250;
// bram[47136] = 253;
// bram[47137] = 253;
// bram[47138] = 248;
// bram[47139] = 241;
// bram[47140] = 229;
// bram[47141] = 215;
// bram[47142] = 198;
// bram[47143] = 179;
// bram[47144] = 158;
// bram[47145] = 136;
// bram[47146] = 115;
// bram[47147] = 93;
// bram[47148] = 72;
// bram[47149] = 53;
// bram[47150] = 37;
// bram[47151] = 23;
// bram[47152] = 12;
// bram[47153] = 4;
// bram[47154] = 0;
// bram[47155] = 0;
// bram[47156] = 3;
// bram[47157] = 11;
// bram[47158] = 21;
// bram[47159] = 35;
// bram[47160] = 52;
// bram[47161] = 71;
// bram[47162] = 91;
// bram[47163] = 113;
// bram[47164] = 134;
// bram[47165] = 156;
// bram[47166] = 177;
// bram[47167] = 196;
// bram[47168] = 213;
// bram[47169] = 228;
// bram[47170] = 240;
// bram[47171] = 248;
// bram[47172] = 252;
// bram[47173] = 253;
// bram[47174] = 250;
// bram[47175] = 244;
// bram[47176] = 234;
// bram[47177] = 220;
// bram[47178] = 204;
// bram[47179] = 186;
// bram[47180] = 166;
// bram[47181] = 144;
// bram[47182] = 123;
// bram[47183] = 101;
// bram[47184] = 80;
// bram[47185] = 60;
// bram[47186] = 43;
// bram[47187] = 27;
// bram[47188] = 15;
// bram[47189] = 6;
// bram[47190] = 1;
// bram[47191] = 0;
// bram[47192] = 2;
// bram[47193] = 8;
// bram[47194] = 17;
// bram[47195] = 30;
// bram[47196] = 46;
// bram[47197] = 64;
// bram[47198] = 83;
// bram[47199] = 105;
// bram[47200] = 127;
// bram[47201] = 148;
// bram[47202] = 170;
// bram[47203] = 189;
// bram[47204] = 207;
// bram[47205] = 223;
// bram[47206] = 236;
// bram[47207] = 245;
// bram[47208] = 251;
// bram[47209] = 253;
// bram[47210] = 252;
// bram[47211] = 247;
// bram[47212] = 238;
// bram[47213] = 226;
// bram[47214] = 210;
// bram[47215] = 193;
// bram[47216] = 173;
// bram[47217] = 152;
// bram[47218] = 130;
// bram[47219] = 109;
// bram[47220] = 87;
// bram[47221] = 67;
// bram[47222] = 49;
// bram[47223] = 33;
// bram[47224] = 19;
// bram[47225] = 9;
// bram[47226] = 3;
// bram[47227] = 0;
// bram[47228] = 1;
// bram[47229] = 5;
// bram[47230] = 13;
// bram[47231] = 25;
// bram[47232] = 40;
// bram[47233] = 57;
// bram[47234] = 76;
// bram[47235] = 97;
// bram[47236] = 119;
// bram[47237] = 140;
// bram[47238] = 162;
// bram[47239] = 182;
// bram[47240] = 201;
// bram[47241] = 218;
// bram[47242] = 232;
// bram[47243] = 242;
// bram[47244] = 250;
// bram[47245] = 253;
// bram[47246] = 253;
// bram[47247] = 249;
// bram[47248] = 241;
// bram[47249] = 230;
// bram[47250] = 216;
// bram[47251] = 200;
// bram[47252] = 181;
// bram[47253] = 160;
// bram[47254] = 138;
// bram[47255] = 117;
// bram[47256] = 95;
// bram[47257] = 74;
// bram[47258] = 55;
// bram[47259] = 38;
// bram[47260] = 24;
// bram[47261] = 12;
// bram[47262] = 5;
// bram[47263] = 0;
// bram[47264] = 0;
// bram[47265] = 3;
// bram[47266] = 10;
// bram[47267] = 20;
// bram[47268] = 34;
// bram[47269] = 50;
// bram[47270] = 69;
// bram[47271] = 89;
// bram[47272] = 111;
// bram[47273] = 132;
// bram[47274] = 154;
// bram[47275] = 175;
// bram[47276] = 195;
// bram[47277] = 212;
// bram[47278] = 227;
// bram[47279] = 239;
// bram[47280] = 247;
// bram[47281] = 252;
// bram[47282] = 253;
// bram[47283] = 251;
// bram[47284] = 245;
// bram[47285] = 235;
// bram[47286] = 222;
// bram[47287] = 206;
// bram[47288] = 188;
// bram[47289] = 168;
// bram[47290] = 146;
// bram[47291] = 125;
// bram[47292] = 103;
// bram[47293] = 82;
// bram[47294] = 62;
// bram[47295] = 44;
// bram[47296] = 29;
// bram[47297] = 16;
// bram[47298] = 7;
// bram[47299] = 1;
// bram[47300] = 0;
// bram[47301] = 1;
// bram[47302] = 7;
// bram[47303] = 16;
// bram[47304] = 29;
// bram[47305] = 44;
// bram[47306] = 62;
// bram[47307] = 82;
// bram[47308] = 103;
// bram[47309] = 125;
// bram[47310] = 146;
// bram[47311] = 168;
// bram[47312] = 188;
// bram[47313] = 206;
// bram[47314] = 222;
// bram[47315] = 235;
// bram[47316] = 245;
// bram[47317] = 251;
// bram[47318] = 253;
// bram[47319] = 252;
// bram[47320] = 247;
// bram[47321] = 239;
// bram[47322] = 227;
// bram[47323] = 212;
// bram[47324] = 195;
// bram[47325] = 175;
// bram[47326] = 154;
// bram[47327] = 132;
// bram[47328] = 111;
// bram[47329] = 89;
// bram[47330] = 69;
// bram[47331] = 50;
// bram[47332] = 34;
// bram[47333] = 20;
// bram[47334] = 10;
// bram[47335] = 3;
// bram[47336] = 0;
// bram[47337] = 0;
// bram[47338] = 5;
// bram[47339] = 12;
// bram[47340] = 24;
// bram[47341] = 38;
// bram[47342] = 55;
// bram[47343] = 74;
// bram[47344] = 95;
// bram[47345] = 117;
// bram[47346] = 138;
// bram[47347] = 160;
// bram[47348] = 181;
// bram[47349] = 200;
// bram[47350] = 216;
// bram[47351] = 230;
// bram[47352] = 241;
// bram[47353] = 249;
// bram[47354] = 253;
// bram[47355] = 253;
// bram[47356] = 250;
// bram[47357] = 242;
// bram[47358] = 232;
// bram[47359] = 218;
// bram[47360] = 201;
// bram[47361] = 182;
// bram[47362] = 162;
// bram[47363] = 140;
// bram[47364] = 119;
// bram[47365] = 97;
// bram[47366] = 76;
// bram[47367] = 57;
// bram[47368] = 40;
// bram[47369] = 25;
// bram[47370] = 13;
// bram[47371] = 5;
// bram[47372] = 1;
// bram[47373] = 0;
// bram[47374] = 3;
// bram[47375] = 9;
// bram[47376] = 19;
// bram[47377] = 33;
// bram[47378] = 49;
// bram[47379] = 67;
// bram[47380] = 87;
// bram[47381] = 109;
// bram[47382] = 130;
// bram[47383] = 152;
// bram[47384] = 173;
// bram[47385] = 193;
// bram[47386] = 210;
// bram[47387] = 226;
// bram[47388] = 238;
// bram[47389] = 247;
// bram[47390] = 252;
// bram[47391] = 253;
// bram[47392] = 251;
// bram[47393] = 245;
// bram[47394] = 236;
// bram[47395] = 223;
// bram[47396] = 207;
// bram[47397] = 189;
// bram[47398] = 170;
// bram[47399] = 148;
// bram[47400] = 126;
// bram[47401] = 105;
// bram[47402] = 83;
// bram[47403] = 64;
// bram[47404] = 46;
// bram[47405] = 30;
// bram[47406] = 17;
// bram[47407] = 8;
// bram[47408] = 2;
// bram[47409] = 0;
// bram[47410] = 1;
// bram[47411] = 6;
// bram[47412] = 15;
// bram[47413] = 27;
// bram[47414] = 43;
// bram[47415] = 60;
// bram[47416] = 80;
// bram[47417] = 101;
// bram[47418] = 123;
// bram[47419] = 144;
// bram[47420] = 166;
// bram[47421] = 186;
// bram[47422] = 204;
// bram[47423] = 220;
// bram[47424] = 234;
// bram[47425] = 244;
// bram[47426] = 250;
// bram[47427] = 253;
// bram[47428] = 252;
// bram[47429] = 248;
// bram[47430] = 240;
// bram[47431] = 228;
// bram[47432] = 213;
// bram[47433] = 196;
// bram[47434] = 177;
// bram[47435] = 156;
// bram[47436] = 134;
// bram[47437] = 113;
// bram[47438] = 91;
// bram[47439] = 71;
// bram[47440] = 52;
// bram[47441] = 35;
// bram[47442] = 21;
// bram[47443] = 11;
// bram[47444] = 3;
// bram[47445] = 0;
// bram[47446] = 0;
// bram[47447] = 4;
// bram[47448] = 12;
// bram[47449] = 23;
// bram[47450] = 37;
// bram[47451] = 53;
// bram[47452] = 72;
// bram[47453] = 93;
// bram[47454] = 115;
// bram[47455] = 136;
// bram[47456] = 158;
// bram[47457] = 179;
// bram[47458] = 198;
// bram[47459] = 215;
// bram[47460] = 229;
// bram[47461] = 241;
// bram[47462] = 248;
// bram[47463] = 253;
// bram[47464] = 253;
// bram[47465] = 250;
// bram[47466] = 243;
// bram[47467] = 233;
// bram[47468] = 219;
// bram[47469] = 203;
// bram[47470] = 184;
// bram[47471] = 164;
// bram[47472] = 142;
// bram[47473] = 121;
// bram[47474] = 99;
// bram[47475] = 78;
// bram[47476] = 58;
// bram[47477] = 41;
// bram[47478] = 26;
// bram[47479] = 14;
// bram[47480] = 6;
// bram[47481] = 1;
// bram[47482] = 0;
// bram[47483] = 2;
// bram[47484] = 8;
// bram[47485] = 18;
// bram[47486] = 31;
// bram[47487] = 47;
// bram[47488] = 65;
// bram[47489] = 85;
// bram[47490] = 107;
// bram[47491] = 128;
// bram[47492] = 150;
// bram[47493] = 171;
// bram[47494] = 191;
// bram[47495] = 209;
// bram[47496] = 224;
// bram[47497] = 237;
// bram[47498] = 246;
// bram[47499] = 252;
// bram[47500] = 254;
// bram[47501] = 252;
// bram[47502] = 246;
// bram[47503] = 237;
// bram[47504] = 224;
// bram[47505] = 209;
// bram[47506] = 191;
// bram[47507] = 171;
// bram[47508] = 150;
// bram[47509] = 128;
// bram[47510] = 107;
// bram[47511] = 85;
// bram[47512] = 65;
// bram[47513] = 47;
// bram[47514] = 31;
// bram[47515] = 18;
// bram[47516] = 8;
// bram[47517] = 2;
// bram[47518] = 0;
// bram[47519] = 1;
// bram[47520] = 6;
// bram[47521] = 14;
// bram[47522] = 26;
// bram[47523] = 41;
// bram[47524] = 58;
// bram[47525] = 78;
// bram[47526] = 99;
// bram[47527] = 121;
// bram[47528] = 142;
// bram[47529] = 164;
// bram[47530] = 184;
// bram[47531] = 203;
// bram[47532] = 219;
// bram[47533] = 233;
// bram[47534] = 243;
// bram[47535] = 250;
// bram[47536] = 253;
// bram[47537] = 253;
// bram[47538] = 248;
// bram[47539] = 241;
// bram[47540] = 229;
// bram[47541] = 215;
// bram[47542] = 198;
// bram[47543] = 179;
// bram[47544] = 158;
// bram[47545] = 136;
// bram[47546] = 115;
// bram[47547] = 93;
// bram[47548] = 72;
// bram[47549] = 53;
// bram[47550] = 37;
// bram[47551] = 23;
// bram[47552] = 12;
// bram[47553] = 4;
// bram[47554] = 0;
// bram[47555] = 0;
// bram[47556] = 3;
// bram[47557] = 11;
// bram[47558] = 21;
// bram[47559] = 35;
// bram[47560] = 52;
// bram[47561] = 71;
// bram[47562] = 91;
// bram[47563] = 113;
// bram[47564] = 134;
// bram[47565] = 156;
// bram[47566] = 177;
// bram[47567] = 196;
// bram[47568] = 213;
// bram[47569] = 228;
// bram[47570] = 240;
// bram[47571] = 248;
// bram[47572] = 252;
// bram[47573] = 253;
// bram[47574] = 250;
// bram[47575] = 244;
// bram[47576] = 234;
// bram[47577] = 220;
// bram[47578] = 204;
// bram[47579] = 186;
// bram[47580] = 166;
// bram[47581] = 144;
// bram[47582] = 123;
// bram[47583] = 101;
// bram[47584] = 80;
// bram[47585] = 60;
// bram[47586] = 43;
// bram[47587] = 27;
// bram[47588] = 15;
// bram[47589] = 6;
// bram[47590] = 1;
// bram[47591] = 0;
// bram[47592] = 2;
// bram[47593] = 8;
// bram[47594] = 17;
// bram[47595] = 30;
// bram[47596] = 46;
// bram[47597] = 64;
// bram[47598] = 83;
// bram[47599] = 105;
// bram[47600] = 127;
// bram[47601] = 148;
// bram[47602] = 170;
// bram[47603] = 189;
// bram[47604] = 207;
// bram[47605] = 223;
// bram[47606] = 236;
// bram[47607] = 245;
// bram[47608] = 251;
// bram[47609] = 253;
// bram[47610] = 252;
// bram[47611] = 247;
// bram[47612] = 238;
// bram[47613] = 226;
// bram[47614] = 210;
// bram[47615] = 193;
// bram[47616] = 173;
// bram[47617] = 152;
// bram[47618] = 130;
// bram[47619] = 109;
// bram[47620] = 87;
// bram[47621] = 67;
// bram[47622] = 49;
// bram[47623] = 33;
// bram[47624] = 19;
// bram[47625] = 9;
// bram[47626] = 3;
// bram[47627] = 0;
// bram[47628] = 1;
// bram[47629] = 5;
// bram[47630] = 13;
// bram[47631] = 25;
// bram[47632] = 40;
// bram[47633] = 57;
// bram[47634] = 76;
// bram[47635] = 97;
// bram[47636] = 119;
// bram[47637] = 140;
// bram[47638] = 162;
// bram[47639] = 182;
// bram[47640] = 201;
// bram[47641] = 218;
// bram[47642] = 232;
// bram[47643] = 242;
// bram[47644] = 250;
// bram[47645] = 253;
// bram[47646] = 253;
// bram[47647] = 249;
// bram[47648] = 241;
// bram[47649] = 230;
// bram[47650] = 216;
// bram[47651] = 200;
// bram[47652] = 181;
// bram[47653] = 160;
// bram[47654] = 138;
// bram[47655] = 117;
// bram[47656] = 95;
// bram[47657] = 74;
// bram[47658] = 55;
// bram[47659] = 38;
// bram[47660] = 24;
// bram[47661] = 12;
// bram[47662] = 5;
// bram[47663] = 0;
// bram[47664] = 0;
// bram[47665] = 3;
// bram[47666] = 10;
// bram[47667] = 20;
// bram[47668] = 34;
// bram[47669] = 50;
// bram[47670] = 69;
// bram[47671] = 89;
// bram[47672] = 111;
// bram[47673] = 132;
// bram[47674] = 154;
// bram[47675] = 175;
// bram[47676] = 195;
// bram[47677] = 212;
// bram[47678] = 227;
// bram[47679] = 239;
// bram[47680] = 247;
// bram[47681] = 252;
// bram[47682] = 253;
// bram[47683] = 251;
// bram[47684] = 245;
// bram[47685] = 235;
// bram[47686] = 222;
// bram[47687] = 206;
// bram[47688] = 188;
// bram[47689] = 168;
// bram[47690] = 146;
// bram[47691] = 125;
// bram[47692] = 103;
// bram[47693] = 82;
// bram[47694] = 62;
// bram[47695] = 44;
// bram[47696] = 29;
// bram[47697] = 16;
// bram[47698] = 7;
// bram[47699] = 1;
// bram[47700] = 0;
// bram[47701] = 1;
// bram[47702] = 7;
// bram[47703] = 16;
// bram[47704] = 29;
// bram[47705] = 44;
// bram[47706] = 62;
// bram[47707] = 82;
// bram[47708] = 103;
// bram[47709] = 125;
// bram[47710] = 146;
// bram[47711] = 168;
// bram[47712] = 188;
// bram[47713] = 206;
// bram[47714] = 222;
// bram[47715] = 235;
// bram[47716] = 245;
// bram[47717] = 251;
// bram[47718] = 253;
// bram[47719] = 252;
// bram[47720] = 247;
// bram[47721] = 239;
// bram[47722] = 227;
// bram[47723] = 212;
// bram[47724] = 195;
// bram[47725] = 175;
// bram[47726] = 154;
// bram[47727] = 132;
// bram[47728] = 111;
// bram[47729] = 89;
// bram[47730] = 69;
// bram[47731] = 50;
// bram[47732] = 34;
// bram[47733] = 20;
// bram[47734] = 10;
// bram[47735] = 3;
// bram[47736] = 0;
// bram[47737] = 0;
// bram[47738] = 5;
// bram[47739] = 12;
// bram[47740] = 24;
// bram[47741] = 38;
// bram[47742] = 55;
// bram[47743] = 74;
// bram[47744] = 95;
// bram[47745] = 117;
// bram[47746] = 138;
// bram[47747] = 160;
// bram[47748] = 181;
// bram[47749] = 200;
// bram[47750] = 216;
// bram[47751] = 230;
// bram[47752] = 241;
// bram[47753] = 249;
// bram[47754] = 253;
// bram[47755] = 253;
// bram[47756] = 250;
// bram[47757] = 242;
// bram[47758] = 232;
// bram[47759] = 218;
// bram[47760] = 201;
// bram[47761] = 182;
// bram[47762] = 162;
// bram[47763] = 140;
// bram[47764] = 119;
// bram[47765] = 97;
// bram[47766] = 76;
// bram[47767] = 57;
// bram[47768] = 40;
// bram[47769] = 25;
// bram[47770] = 13;
// bram[47771] = 5;
// bram[47772] = 1;
// bram[47773] = 0;
// bram[47774] = 3;
// bram[47775] = 9;
// bram[47776] = 19;
// bram[47777] = 33;
// bram[47778] = 49;
// bram[47779] = 67;
// bram[47780] = 87;
// bram[47781] = 109;
// bram[47782] = 130;
// bram[47783] = 152;
// bram[47784] = 173;
// bram[47785] = 193;
// bram[47786] = 210;
// bram[47787] = 226;
// bram[47788] = 238;
// bram[47789] = 247;
// bram[47790] = 252;
// bram[47791] = 253;
// bram[47792] = 251;
// bram[47793] = 245;
// bram[47794] = 236;
// bram[47795] = 223;
// bram[47796] = 207;
// bram[47797] = 189;
// bram[47798] = 170;
// bram[47799] = 148;
// bram[47800] = 126;
// bram[47801] = 105;
// bram[47802] = 83;
// bram[47803] = 64;
// bram[47804] = 46;
// bram[47805] = 30;
// bram[47806] = 17;
// bram[47807] = 8;
// bram[47808] = 2;
// bram[47809] = 0;
// bram[47810] = 1;
// bram[47811] = 6;
// bram[47812] = 15;
// bram[47813] = 27;
// bram[47814] = 43;
// bram[47815] = 60;
// bram[47816] = 80;
// bram[47817] = 101;
// bram[47818] = 123;
// bram[47819] = 144;
// bram[47820] = 166;
// bram[47821] = 186;
// bram[47822] = 204;
// bram[47823] = 220;
// bram[47824] = 234;
// bram[47825] = 244;
// bram[47826] = 250;
// bram[47827] = 253;
// bram[47828] = 252;
// bram[47829] = 248;
// bram[47830] = 240;
// bram[47831] = 228;
// bram[47832] = 213;
// bram[47833] = 196;
// bram[47834] = 177;
// bram[47835] = 156;
// bram[47836] = 134;
// bram[47837] = 113;
// bram[47838] = 91;
// bram[47839] = 71;
// bram[47840] = 52;
// bram[47841] = 35;
// bram[47842] = 21;
// bram[47843] = 11;
// bram[47844] = 3;
// bram[47845] = 0;
// bram[47846] = 0;
// bram[47847] = 4;
// bram[47848] = 12;
// bram[47849] = 23;
// bram[47850] = 37;
// bram[47851] = 53;
// bram[47852] = 72;
// bram[47853] = 93;
// bram[47854] = 115;
// bram[47855] = 136;
// bram[47856] = 158;
// bram[47857] = 179;
// bram[47858] = 198;
// bram[47859] = 215;
// bram[47860] = 229;
// bram[47861] = 241;
// bram[47862] = 248;
// bram[47863] = 253;
// bram[47864] = 253;
// bram[47865] = 250;
// bram[47866] = 243;
// bram[47867] = 233;
// bram[47868] = 219;
// bram[47869] = 203;
// bram[47870] = 184;
// bram[47871] = 164;
// bram[47872] = 142;
// bram[47873] = 121;
// bram[47874] = 99;
// bram[47875] = 78;
// bram[47876] = 58;
// bram[47877] = 41;
// bram[47878] = 26;
// bram[47879] = 14;
// bram[47880] = 6;
// bram[47881] = 1;
// bram[47882] = 0;
// bram[47883] = 2;
// bram[47884] = 8;
// bram[47885] = 18;
// bram[47886] = 31;
// bram[47887] = 47;
// bram[47888] = 65;
// bram[47889] = 85;
// bram[47890] = 107;
// bram[47891] = 128;
// bram[47892] = 150;
// bram[47893] = 171;
// bram[47894] = 191;
// bram[47895] = 209;
// bram[47896] = 224;
// bram[47897] = 237;
// bram[47898] = 246;
// bram[47899] = 252;
// bram[47900] = 254;
// bram[47901] = 252;
// bram[47902] = 246;
// bram[47903] = 237;
// bram[47904] = 224;
// bram[47905] = 209;
// bram[47906] = 191;
// bram[47907] = 171;
// bram[47908] = 150;
// bram[47909] = 128;
// bram[47910] = 107;
// bram[47911] = 85;
// bram[47912] = 65;
// bram[47913] = 47;
// bram[47914] = 31;
// bram[47915] = 18;
// bram[47916] = 8;
// bram[47917] = 2;
// bram[47918] = 0;
// bram[47919] = 1;
// bram[47920] = 6;
// bram[47921] = 14;
// bram[47922] = 26;
// bram[47923] = 41;
// bram[47924] = 58;
// bram[47925] = 78;
// bram[47926] = 99;
// bram[47927] = 121;
// bram[47928] = 142;
// bram[47929] = 164;
// bram[47930] = 184;
// bram[47931] = 203;
// bram[47932] = 219;
// bram[47933] = 233;
// bram[47934] = 243;
// bram[47935] = 250;
// bram[47936] = 253;
// bram[47937] = 253;
// bram[47938] = 248;
// bram[47939] = 241;
// bram[47940] = 229;
// bram[47941] = 215;
// bram[47942] = 198;
// bram[47943] = 179;
// bram[47944] = 158;
// bram[47945] = 136;
// bram[47946] = 115;
// bram[47947] = 93;
// bram[47948] = 72;
// bram[47949] = 53;
// bram[47950] = 37;
// bram[47951] = 23;
// bram[47952] = 12;
// bram[47953] = 4;
// bram[47954] = 0;
// bram[47955] = 0;
// bram[47956] = 3;
// bram[47957] = 11;
// bram[47958] = 21;
// bram[47959] = 35;
// bram[47960] = 52;
// bram[47961] = 71;
// bram[47962] = 91;
// bram[47963] = 113;
// bram[47964] = 134;
// bram[47965] = 156;
// bram[47966] = 177;
// bram[47967] = 196;
// bram[47968] = 213;
// bram[47969] = 228;
// bram[47970] = 240;
// bram[47971] = 248;
// bram[47972] = 252;
// bram[47973] = 253;
// bram[47974] = 250;
// bram[47975] = 244;
// bram[47976] = 234;
// bram[47977] = 220;
// bram[47978] = 204;
// bram[47979] = 186;
// bram[47980] = 166;
// bram[47981] = 144;
// bram[47982] = 123;
// bram[47983] = 101;
// bram[47984] = 80;
// bram[47985] = 60;
// bram[47986] = 43;
// bram[47987] = 27;
// bram[47988] = 15;
// bram[47989] = 6;
// bram[47990] = 1;
// bram[47991] = 0;
// bram[47992] = 2;
// bram[47993] = 8;
// bram[47994] = 17;
// bram[47995] = 30;
// bram[47996] = 46;
// bram[47997] = 64;
// bram[47998] = 83;
// bram[47999] = 105;
// bram[48000] = 127;
// bram[48001] = 151;
// bram[48002] = 174;
// bram[48003] = 196;
// bram[48004] = 215;
// bram[48005] = 231;
// bram[48006] = 243;
// bram[48007] = 251;
// bram[48008] = 253;
// bram[48009] = 252;
// bram[48010] = 245;
// bram[48011] = 234;
// bram[48012] = 219;
// bram[48013] = 201;
// bram[48014] = 180;
// bram[48015] = 156;
// bram[48016] = 132;
// bram[48017] = 108;
// bram[48018] = 84;
// bram[48019] = 62;
// bram[48020] = 42;
// bram[48021] = 25;
// bram[48022] = 12;
// bram[48023] = 4;
// bram[48024] = 0;
// bram[48025] = 1;
// bram[48026] = 6;
// bram[48027] = 16;
// bram[48028] = 30;
// bram[48029] = 48;
// bram[48030] = 68;
// bram[48031] = 91;
// bram[48032] = 115;
// bram[48033] = 140;
// bram[48034] = 164;
// bram[48035] = 187;
// bram[48036] = 207;
// bram[48037] = 224;
// bram[48038] = 238;
// bram[48039] = 248;
// bram[48040] = 253;
// bram[48041] = 253;
// bram[48042] = 249;
// bram[48043] = 240;
// bram[48044] = 226;
// bram[48045] = 210;
// bram[48046] = 190;
// bram[48047] = 167;
// bram[48048] = 143;
// bram[48049] = 119;
// bram[48050] = 94;
// bram[48051] = 71;
// bram[48052] = 50;
// bram[48053] = 32;
// bram[48054] = 18;
// bram[48055] = 7;
// bram[48056] = 1;
// bram[48057] = 0;
// bram[48058] = 3;
// bram[48059] = 11;
// bram[48060] = 23;
// bram[48061] = 39;
// bram[48062] = 59;
// bram[48063] = 81;
// bram[48064] = 104;
// bram[48065] = 129;
// bram[48066] = 153;
// bram[48067] = 177;
// bram[48068] = 198;
// bram[48069] = 217;
// bram[48070] = 232;
// bram[48071] = 244;
// bram[48072] = 251;
// bram[48073] = 253;
// bram[48074] = 251;
// bram[48075] = 244;
// bram[48076] = 233;
// bram[48077] = 218;
// bram[48078] = 199;
// bram[48079] = 178;
// bram[48080] = 154;
// bram[48081] = 130;
// bram[48082] = 105;
// bram[48083] = 82;
// bram[48084] = 60;
// bram[48085] = 40;
// bram[48086] = 24;
// bram[48087] = 11;
// bram[48088] = 3;
// bram[48089] = 0;
// bram[48090] = 1;
// bram[48091] = 7;
// bram[48092] = 17;
// bram[48093] = 32;
// bram[48094] = 50;
// bram[48095] = 70;
// bram[48096] = 93;
// bram[48097] = 118;
// bram[48098] = 142;
// bram[48099] = 166;
// bram[48100] = 189;
// bram[48101] = 209;
// bram[48102] = 226;
// bram[48103] = 239;
// bram[48104] = 248;
// bram[48105] = 253;
// bram[48106] = 253;
// bram[48107] = 248;
// bram[48108] = 239;
// bram[48109] = 225;
// bram[48110] = 208;
// bram[48111] = 188;
// bram[48112] = 165;
// bram[48113] = 141;
// bram[48114] = 116;
// bram[48115] = 92;
// bram[48116] = 69;
// bram[48117] = 49;
// bram[48118] = 31;
// bram[48119] = 17;
// bram[48120] = 6;
// bram[48121] = 1;
// bram[48122] = 0;
// bram[48123] = 3;
// bram[48124] = 12;
// bram[48125] = 24;
// bram[48126] = 41;
// bram[48127] = 61;
// bram[48128] = 83;
// bram[48129] = 106;
// bram[48130] = 131;
// bram[48131] = 155;
// bram[48132] = 179;
// bram[48133] = 200;
// bram[48134] = 218;
// bram[48135] = 234;
// bram[48136] = 245;
// bram[48137] = 251;
// bram[48138] = 253;
// bram[48139] = 251;
// bram[48140] = 243;
// bram[48141] = 232;
// bram[48142] = 216;
// bram[48143] = 197;
// bram[48144] = 175;
// bram[48145] = 152;
// bram[48146] = 128;
// bram[48147] = 103;
// bram[48148] = 80;
// bram[48149] = 58;
// bram[48150] = 38;
// bram[48151] = 23;
// bram[48152] = 10;
// bram[48153] = 3;
// bram[48154] = 0;
// bram[48155] = 1;
// bram[48156] = 7;
// bram[48157] = 18;
// bram[48158] = 33;
// bram[48159] = 51;
// bram[48160] = 72;
// bram[48161] = 96;
// bram[48162] = 120;
// bram[48163] = 144;
// bram[48164] = 168;
// bram[48165] = 191;
// bram[48166] = 210;
// bram[48167] = 227;
// bram[48168] = 240;
// bram[48169] = 249;
// bram[48170] = 253;
// bram[48171] = 253;
// bram[48172] = 247;
// bram[48173] = 238;
// bram[48174] = 224;
// bram[48175] = 206;
// bram[48176] = 186;
// bram[48177] = 163;
// bram[48178] = 139;
// bram[48179] = 114;
// bram[48180] = 90;
// bram[48181] = 67;
// bram[48182] = 47;
// bram[48183] = 29;
// bram[48184] = 15;
// bram[48185] = 6;
// bram[48186] = 0;
// bram[48187] = 0;
// bram[48188] = 4;
// bram[48189] = 13;
// bram[48190] = 26;
// bram[48191] = 43;
// bram[48192] = 63;
// bram[48193] = 85;
// bram[48194] = 109;
// bram[48195] = 133;
// bram[48196] = 158;
// bram[48197] = 181;
// bram[48198] = 202;
// bram[48199] = 220;
// bram[48200] = 235;
// bram[48201] = 246;
// bram[48202] = 252;
// bram[48203] = 253;
// bram[48204] = 250;
// bram[48205] = 243;
// bram[48206] = 230;
// bram[48207] = 214;
// bram[48208] = 195;
// bram[48209] = 173;
// bram[48210] = 150;
// bram[48211] = 125;
// bram[48212] = 101;
// bram[48213] = 77;
// bram[48214] = 56;
// bram[48215] = 37;
// bram[48216] = 21;
// bram[48217] = 10;
// bram[48218] = 2;
// bram[48219] = 0;
// bram[48220] = 2;
// bram[48221] = 8;
// bram[48222] = 19;
// bram[48223] = 35;
// bram[48224] = 53;
// bram[48225] = 74;
// bram[48226] = 98;
// bram[48227] = 122;
// bram[48228] = 147;
// bram[48229] = 170;
// bram[48230] = 192;
// bram[48231] = 212;
// bram[48232] = 229;
// bram[48233] = 241;
// bram[48234] = 250;
// bram[48235] = 253;
// bram[48236] = 252;
// bram[48237] = 247;
// bram[48238] = 236;
// bram[48239] = 222;
// bram[48240] = 204;
// bram[48241] = 184;
// bram[48242] = 161;
// bram[48243] = 137;
// bram[48244] = 112;
// bram[48245] = 88;
// bram[48246] = 65;
// bram[48247] = 45;
// bram[48248] = 28;
// bram[48249] = 14;
// bram[48250] = 5;
// bram[48251] = 0;
// bram[48252] = 0;
// bram[48253] = 5;
// bram[48254] = 14;
// bram[48255] = 27;
// bram[48256] = 44;
// bram[48257] = 64;
// bram[48258] = 87;
// bram[48259] = 111;
// bram[48260] = 135;
// bram[48261] = 160;
// bram[48262] = 183;
// bram[48263] = 204;
// bram[48264] = 221;
// bram[48265] = 236;
// bram[48266] = 246;
// bram[48267] = 252;
// bram[48268] = 253;
// bram[48269] = 250;
// bram[48270] = 242;
// bram[48271] = 229;
// bram[48272] = 213;
// bram[48273] = 193;
// bram[48274] = 171;
// bram[48275] = 148;
// bram[48276] = 123;
// bram[48277] = 99;
// bram[48278] = 75;
// bram[48279] = 54;
// bram[48280] = 35;
// bram[48281] = 20;
// bram[48282] = 9;
// bram[48283] = 2;
// bram[48284] = 0;
// bram[48285] = 2;
// bram[48286] = 9;
// bram[48287] = 21;
// bram[48288] = 36;
// bram[48289] = 55;
// bram[48290] = 77;
// bram[48291] = 100;
// bram[48292] = 124;
// bram[48293] = 149;
// bram[48294] = 172;
// bram[48295] = 194;
// bram[48296] = 214;
// bram[48297] = 230;
// bram[48298] = 242;
// bram[48299] = 250;
// bram[48300] = 253;
// bram[48301] = 252;
// bram[48302] = 246;
// bram[48303] = 235;
// bram[48304] = 221;
// bram[48305] = 203;
// bram[48306] = 182;
// bram[48307] = 159;
// bram[48308] = 134;
// bram[48309] = 110;
// bram[48310] = 86;
// bram[48311] = 63;
// bram[48312] = 43;
// bram[48313] = 26;
// bram[48314] = 13;
// bram[48315] = 4;
// bram[48316] = 0;
// bram[48317] = 0;
// bram[48318] = 5;
// bram[48319] = 15;
// bram[48320] = 29;
// bram[48321] = 46;
// bram[48322] = 66;
// bram[48323] = 89;
// bram[48324] = 113;
// bram[48325] = 138;
// bram[48326] = 162;
// bram[48327] = 185;
// bram[48328] = 205;
// bram[48329] = 223;
// bram[48330] = 237;
// bram[48331] = 247;
// bram[48332] = 252;
// bram[48333] = 253;
// bram[48334] = 249;
// bram[48335] = 241;
// bram[48336] = 228;
// bram[48337] = 211;
// bram[48338] = 191;
// bram[48339] = 169;
// bram[48340] = 145;
// bram[48341] = 121;
// bram[48342] = 97;
// bram[48343] = 73;
// bram[48344] = 52;
// bram[48345] = 34;
// bram[48346] = 19;
// bram[48347] = 8;
// bram[48348] = 1;
// bram[48349] = 0;
// bram[48350] = 2;
// bram[48351] = 10;
// bram[48352] = 22;
// bram[48353] = 38;
// bram[48354] = 57;
// bram[48355] = 79;
// bram[48356] = 102;
// bram[48357] = 127;
// bram[48358] = 151;
// bram[48359] = 175;
// bram[48360] = 196;
// bram[48361] = 215;
// bram[48362] = 231;
// bram[48363] = 243;
// bram[48364] = 251;
// bram[48365] = 253;
// bram[48366] = 252;
// bram[48367] = 245;
// bram[48368] = 234;
// bram[48369] = 219;
// bram[48370] = 201;
// bram[48371] = 180;
// bram[48372] = 156;
// bram[48373] = 132;
// bram[48374] = 108;
// bram[48375] = 84;
// bram[48376] = 62;
// bram[48377] = 42;
// bram[48378] = 25;
// bram[48379] = 12;
// bram[48380] = 4;
// bram[48381] = 0;
// bram[48382] = 1;
// bram[48383] = 6;
// bram[48384] = 16;
// bram[48385] = 30;
// bram[48386] = 48;
// bram[48387] = 68;
// bram[48388] = 91;
// bram[48389] = 115;
// bram[48390] = 140;
// bram[48391] = 164;
// bram[48392] = 187;
// bram[48393] = 207;
// bram[48394] = 224;
// bram[48395] = 238;
// bram[48396] = 248;
// bram[48397] = 253;
// bram[48398] = 253;
// bram[48399] = 249;
// bram[48400] = 240;
// bram[48401] = 226;
// bram[48402] = 210;
// bram[48403] = 189;
// bram[48404] = 167;
// bram[48405] = 143;
// bram[48406] = 119;
// bram[48407] = 94;
// bram[48408] = 71;
// bram[48409] = 50;
// bram[48410] = 32;
// bram[48411] = 18;
// bram[48412] = 7;
// bram[48413] = 1;
// bram[48414] = 0;
// bram[48415] = 3;
// bram[48416] = 11;
// bram[48417] = 23;
// bram[48418] = 39;
// bram[48419] = 59;
// bram[48420] = 81;
// bram[48421] = 104;
// bram[48422] = 129;
// bram[48423] = 153;
// bram[48424] = 177;
// bram[48425] = 198;
// bram[48426] = 217;
// bram[48427] = 232;
// bram[48428] = 244;
// bram[48429] = 251;
// bram[48430] = 253;
// bram[48431] = 251;
// bram[48432] = 244;
// bram[48433] = 233;
// bram[48434] = 218;
// bram[48435] = 199;
// bram[48436] = 177;
// bram[48437] = 154;
// bram[48438] = 130;
// bram[48439] = 105;
// bram[48440] = 82;
// bram[48441] = 60;
// bram[48442] = 40;
// bram[48443] = 24;
// bram[48444] = 11;
// bram[48445] = 3;
// bram[48446] = 0;
// bram[48447] = 1;
// bram[48448] = 7;
// bram[48449] = 17;
// bram[48450] = 32;
// bram[48451] = 50;
// bram[48452] = 70;
// bram[48453] = 93;
// bram[48454] = 118;
// bram[48455] = 142;
// bram[48456] = 166;
// bram[48457] = 189;
// bram[48458] = 209;
// bram[48459] = 226;
// bram[48460] = 239;
// bram[48461] = 248;
// bram[48462] = 253;
// bram[48463] = 253;
// bram[48464] = 248;
// bram[48465] = 239;
// bram[48466] = 225;
// bram[48467] = 208;
// bram[48468] = 188;
// bram[48469] = 165;
// bram[48470] = 141;
// bram[48471] = 116;
// bram[48472] = 92;
// bram[48473] = 69;
// bram[48474] = 49;
// bram[48475] = 31;
// bram[48476] = 16;
// bram[48477] = 6;
// bram[48478] = 1;
// bram[48479] = 0;
// bram[48480] = 3;
// bram[48481] = 12;
// bram[48482] = 25;
// bram[48483] = 41;
// bram[48484] = 61;
// bram[48485] = 83;
// bram[48486] = 107;
// bram[48487] = 131;
// bram[48488] = 155;
// bram[48489] = 179;
// bram[48490] = 200;
// bram[48491] = 218;
// bram[48492] = 234;
// bram[48493] = 245;
// bram[48494] = 251;
// bram[48495] = 253;
// bram[48496] = 251;
// bram[48497] = 243;
// bram[48498] = 232;
// bram[48499] = 216;
// bram[48500] = 197;
// bram[48501] = 175;
// bram[48502] = 152;
// bram[48503] = 128;
// bram[48504] = 103;
// bram[48505] = 80;
// bram[48506] = 58;
// bram[48507] = 38;
// bram[48508] = 22;
// bram[48509] = 10;
// bram[48510] = 3;
// bram[48511] = 0;
// bram[48512] = 1;
// bram[48513] = 8;
// bram[48514] = 18;
// bram[48515] = 33;
// bram[48516] = 51;
// bram[48517] = 72;
// bram[48518] = 96;
// bram[48519] = 120;
// bram[48520] = 144;
// bram[48521] = 168;
// bram[48522] = 191;
// bram[48523] = 210;
// bram[48524] = 227;
// bram[48525] = 240;
// bram[48526] = 249;
// bram[48527] = 253;
// bram[48528] = 253;
// bram[48529] = 247;
// bram[48530] = 238;
// bram[48531] = 224;
// bram[48532] = 206;
// bram[48533] = 186;
// bram[48534] = 163;
// bram[48535] = 139;
// bram[48536] = 114;
// bram[48537] = 90;
// bram[48538] = 67;
// bram[48539] = 47;
// bram[48540] = 29;
// bram[48541] = 15;
// bram[48542] = 6;
// bram[48543] = 0;
// bram[48544] = 0;
// bram[48545] = 4;
// bram[48546] = 13;
// bram[48547] = 26;
// bram[48548] = 43;
// bram[48549] = 63;
// bram[48550] = 85;
// bram[48551] = 109;
// bram[48552] = 133;
// bram[48553] = 158;
// bram[48554] = 181;
// bram[48555] = 202;
// bram[48556] = 220;
// bram[48557] = 235;
// bram[48558] = 246;
// bram[48559] = 252;
// bram[48560] = 253;
// bram[48561] = 250;
// bram[48562] = 243;
// bram[48563] = 230;
// bram[48564] = 214;
// bram[48565] = 195;
// bram[48566] = 173;
// bram[48567] = 150;
// bram[48568] = 125;
// bram[48569] = 101;
// bram[48570] = 77;
// bram[48571] = 56;
// bram[48572] = 37;
// bram[48573] = 21;
// bram[48574] = 10;
// bram[48575] = 2;
// bram[48576] = 0;
// bram[48577] = 2;
// bram[48578] = 8;
// bram[48579] = 19;
// bram[48580] = 35;
// bram[48581] = 53;
// bram[48582] = 75;
// bram[48583] = 98;
// bram[48584] = 122;
// bram[48585] = 147;
// bram[48586] = 170;
// bram[48587] = 192;
// bram[48588] = 212;
// bram[48589] = 229;
// bram[48590] = 241;
// bram[48591] = 250;
// bram[48592] = 253;
// bram[48593] = 252;
// bram[48594] = 247;
// bram[48595] = 236;
// bram[48596] = 222;
// bram[48597] = 204;
// bram[48598] = 184;
// bram[48599] = 161;
// bram[48600] = 136;
// bram[48601] = 112;
// bram[48602] = 88;
// bram[48603] = 65;
// bram[48604] = 45;
// bram[48605] = 28;
// bram[48606] = 14;
// bram[48607] = 5;
// bram[48608] = 0;
// bram[48609] = 0;
// bram[48610] = 5;
// bram[48611] = 14;
// bram[48612] = 27;
// bram[48613] = 44;
// bram[48614] = 65;
// bram[48615] = 87;
// bram[48616] = 111;
// bram[48617] = 136;
// bram[48618] = 160;
// bram[48619] = 183;
// bram[48620] = 204;
// bram[48621] = 222;
// bram[48622] = 236;
// bram[48623] = 246;
// bram[48624] = 252;
// bram[48625] = 253;
// bram[48626] = 250;
// bram[48627] = 242;
// bram[48628] = 229;
// bram[48629] = 213;
// bram[48630] = 193;
// bram[48631] = 171;
// bram[48632] = 148;
// bram[48633] = 123;
// bram[48634] = 99;
// bram[48635] = 75;
// bram[48636] = 54;
// bram[48637] = 35;
// bram[48638] = 20;
// bram[48639] = 9;
// bram[48640] = 2;
// bram[48641] = 0;
// bram[48642] = 2;
// bram[48643] = 9;
// bram[48644] = 21;
// bram[48645] = 36;
// bram[48646] = 55;
// bram[48647] = 77;
// bram[48648] = 100;
// bram[48649] = 124;
// bram[48650] = 149;
// bram[48651] = 172;
// bram[48652] = 194;
// bram[48653] = 214;
// bram[48654] = 230;
// bram[48655] = 242;
// bram[48656] = 250;
// bram[48657] = 253;
// bram[48658] = 252;
// bram[48659] = 246;
// bram[48660] = 235;
// bram[48661] = 221;
// bram[48662] = 203;
// bram[48663] = 182;
// bram[48664] = 158;
// bram[48665] = 134;
// bram[48666] = 110;
// bram[48667] = 86;
// bram[48668] = 63;
// bram[48669] = 43;
// bram[48670] = 26;
// bram[48671] = 13;
// bram[48672] = 4;
// bram[48673] = 0;
// bram[48674] = 0;
// bram[48675] = 5;
// bram[48676] = 15;
// bram[48677] = 29;
// bram[48678] = 46;
// bram[48679] = 67;
// bram[48680] = 89;
// bram[48681] = 113;
// bram[48682] = 138;
// bram[48683] = 162;
// bram[48684] = 185;
// bram[48685] = 205;
// bram[48686] = 223;
// bram[48687] = 237;
// bram[48688] = 247;
// bram[48689] = 252;
// bram[48690] = 253;
// bram[48691] = 249;
// bram[48692] = 241;
// bram[48693] = 228;
// bram[48694] = 211;
// bram[48695] = 191;
// bram[48696] = 169;
// bram[48697] = 145;
// bram[48698] = 121;
// bram[48699] = 97;
// bram[48700] = 73;
// bram[48701] = 52;
// bram[48702] = 34;
// bram[48703] = 19;
// bram[48704] = 8;
// bram[48705] = 1;
// bram[48706] = 0;
// bram[48707] = 2;
// bram[48708] = 10;
// bram[48709] = 22;
// bram[48710] = 38;
// bram[48711] = 57;
// bram[48712] = 79;
// bram[48713] = 102;
// bram[48714] = 127;
// bram[48715] = 151;
// bram[48716] = 175;
// bram[48717] = 196;
// bram[48718] = 215;
// bram[48719] = 231;
// bram[48720] = 243;
// bram[48721] = 251;
// bram[48722] = 253;
// bram[48723] = 252;
// bram[48724] = 245;
// bram[48725] = 234;
// bram[48726] = 219;
// bram[48727] = 201;
// bram[48728] = 179;
// bram[48729] = 156;
// bram[48730] = 132;
// bram[48731] = 107;
// bram[48732] = 84;
// bram[48733] = 61;
// bram[48734] = 42;
// bram[48735] = 25;
// bram[48736] = 12;
// bram[48737] = 4;
// bram[48738] = 0;
// bram[48739] = 1;
// bram[48740] = 6;
// bram[48741] = 16;
// bram[48742] = 30;
// bram[48743] = 48;
// bram[48744] = 68;
// bram[48745] = 91;
// bram[48746] = 115;
// bram[48747] = 140;
// bram[48748] = 164;
// bram[48749] = 187;
// bram[48750] = 207;
// bram[48751] = 224;
// bram[48752] = 238;
// bram[48753] = 248;
// bram[48754] = 253;
// bram[48755] = 253;
// bram[48756] = 249;
// bram[48757] = 240;
// bram[48758] = 226;
// bram[48759] = 209;
// bram[48760] = 189;
// bram[48761] = 167;
// bram[48762] = 143;
// bram[48763] = 119;
// bram[48764] = 94;
// bram[48765] = 71;
// bram[48766] = 50;
// bram[48767] = 32;
// bram[48768] = 18;
// bram[48769] = 7;
// bram[48770] = 1;
// bram[48771] = 0;
// bram[48772] = 3;
// bram[48773] = 11;
// bram[48774] = 23;
// bram[48775] = 39;
// bram[48776] = 59;
// bram[48777] = 81;
// bram[48778] = 104;
// bram[48779] = 129;
// bram[48780] = 153;
// bram[48781] = 177;
// bram[48782] = 198;
// bram[48783] = 217;
// bram[48784] = 232;
// bram[48785] = 244;
// bram[48786] = 251;
// bram[48787] = 253;
// bram[48788] = 251;
// bram[48789] = 244;
// bram[48790] = 233;
// bram[48791] = 218;
// bram[48792] = 199;
// bram[48793] = 177;
// bram[48794] = 154;
// bram[48795] = 130;
// bram[48796] = 105;
// bram[48797] = 82;
// bram[48798] = 60;
// bram[48799] = 40;
// bram[48800] = 24;
// bram[48801] = 11;
// bram[48802] = 3;
// bram[48803] = 0;
// bram[48804] = 1;
// bram[48805] = 7;
// bram[48806] = 17;
// bram[48807] = 32;
// bram[48808] = 50;
// bram[48809] = 70;
// bram[48810] = 93;
// bram[48811] = 118;
// bram[48812] = 142;
// bram[48813] = 166;
// bram[48814] = 189;
// bram[48815] = 209;
// bram[48816] = 226;
// bram[48817] = 239;
// bram[48818] = 248;
// bram[48819] = 253;
// bram[48820] = 253;
// bram[48821] = 248;
// bram[48822] = 239;
// bram[48823] = 225;
// bram[48824] = 208;
// bram[48825] = 187;
// bram[48826] = 165;
// bram[48827] = 141;
// bram[48828] = 116;
// bram[48829] = 92;
// bram[48830] = 69;
// bram[48831] = 49;
// bram[48832] = 31;
// bram[48833] = 16;
// bram[48834] = 6;
// bram[48835] = 1;
// bram[48836] = 0;
// bram[48837] = 4;
// bram[48838] = 12;
// bram[48839] = 25;
// bram[48840] = 41;
// bram[48841] = 61;
// bram[48842] = 83;
// bram[48843] = 107;
// bram[48844] = 131;
// bram[48845] = 155;
// bram[48846] = 179;
// bram[48847] = 200;
// bram[48848] = 219;
// bram[48849] = 234;
// bram[48850] = 245;
// bram[48851] = 251;
// bram[48852] = 253;
// bram[48853] = 251;
// bram[48854] = 243;
// bram[48855] = 232;
// bram[48856] = 216;
// bram[48857] = 197;
// bram[48858] = 175;
// bram[48859] = 152;
// bram[48860] = 127;
// bram[48861] = 103;
// bram[48862] = 79;
// bram[48863] = 58;
// bram[48864] = 38;
// bram[48865] = 22;
// bram[48866] = 10;
// bram[48867] = 3;
// bram[48868] = 0;
// bram[48869] = 1;
// bram[48870] = 8;
// bram[48871] = 18;
// bram[48872] = 33;
// bram[48873] = 51;
// bram[48874] = 73;
// bram[48875] = 96;
// bram[48876] = 120;
// bram[48877] = 144;
// bram[48878] = 168;
// bram[48879] = 191;
// bram[48880] = 210;
// bram[48881] = 227;
// bram[48882] = 240;
// bram[48883] = 249;
// bram[48884] = 253;
// bram[48885] = 253;
// bram[48886] = 247;
// bram[48887] = 238;
// bram[48888] = 224;
// bram[48889] = 206;
// bram[48890] = 185;
// bram[48891] = 163;
// bram[48892] = 139;
// bram[48893] = 114;
// bram[48894] = 90;
// bram[48895] = 67;
// bram[48896] = 47;
// bram[48897] = 29;
// bram[48898] = 15;
// bram[48899] = 6;
// bram[48900] = 0;
// bram[48901] = 0;
// bram[48902] = 4;
// bram[48903] = 13;
// bram[48904] = 26;
// bram[48905] = 43;
// bram[48906] = 63;
// bram[48907] = 85;
// bram[48908] = 109;
// bram[48909] = 133;
// bram[48910] = 158;
// bram[48911] = 181;
// bram[48912] = 202;
// bram[48913] = 220;
// bram[48914] = 235;
// bram[48915] = 246;
// bram[48916] = 252;
// bram[48917] = 253;
// bram[48918] = 250;
// bram[48919] = 243;
// bram[48920] = 230;
// bram[48921] = 214;
// bram[48922] = 195;
// bram[48923] = 173;
// bram[48924] = 150;
// bram[48925] = 125;
// bram[48926] = 101;
// bram[48927] = 77;
// bram[48928] = 56;
// bram[48929] = 37;
// bram[48930] = 21;
// bram[48931] = 9;
// bram[48932] = 2;
// bram[48933] = 0;
// bram[48934] = 2;
// bram[48935] = 8;
// bram[48936] = 19;
// bram[48937] = 35;
// bram[48938] = 53;
// bram[48939] = 75;
// bram[48940] = 98;
// bram[48941] = 122;
// bram[48942] = 147;
// bram[48943] = 170;
// bram[48944] = 193;
// bram[48945] = 212;
// bram[48946] = 229;
// bram[48947] = 241;
// bram[48948] = 250;
// bram[48949] = 253;
// bram[48950] = 252;
// bram[48951] = 247;
// bram[48952] = 236;
// bram[48953] = 222;
// bram[48954] = 204;
// bram[48955] = 183;
// bram[48956] = 161;
// bram[48957] = 136;
// bram[48958] = 112;
// bram[48959] = 88;
// bram[48960] = 65;
// bram[48961] = 45;
// bram[48962] = 28;
// bram[48963] = 14;
// bram[48964] = 5;
// bram[48965] = 0;
// bram[48966] = 0;
// bram[48967] = 5;
// bram[48968] = 14;
// bram[48969] = 27;
// bram[48970] = 44;
// bram[48971] = 65;
// bram[48972] = 87;
// bram[48973] = 111;
// bram[48974] = 136;
// bram[48975] = 160;
// bram[48976] = 183;
// bram[48977] = 204;
// bram[48978] = 222;
// bram[48979] = 236;
// bram[48980] = 246;
// bram[48981] = 252;
// bram[48982] = 253;
// bram[48983] = 250;
// bram[48984] = 242;
// bram[48985] = 229;
// bram[48986] = 213;
// bram[48987] = 193;
// bram[48988] = 171;
// bram[48989] = 147;
// bram[48990] = 123;
// bram[48991] = 99;
// bram[48992] = 75;
// bram[48993] = 54;
// bram[48994] = 35;
// bram[48995] = 20;
// bram[48996] = 9;
// bram[48997] = 2;
// bram[48998] = 0;
// bram[48999] = 2;
// bram[49000] = 9;
// bram[49001] = 21;
// bram[49002] = 36;
// bram[49003] = 55;
// bram[49004] = 77;
// bram[49005] = 100;
// bram[49006] = 124;
// bram[49007] = 149;
// bram[49008] = 173;
// bram[49009] = 194;
// bram[49010] = 214;
// bram[49011] = 230;
// bram[49012] = 242;
// bram[49013] = 250;
// bram[49014] = 253;
// bram[49015] = 252;
// bram[49016] = 246;
// bram[49017] = 235;
// bram[49018] = 221;
// bram[49019] = 202;
// bram[49020] = 181;
// bram[49021] = 158;
// bram[49022] = 134;
// bram[49023] = 110;
// bram[49024] = 86;
// bram[49025] = 63;
// bram[49026] = 43;
// bram[49027] = 26;
// bram[49028] = 13;
// bram[49029] = 4;
// bram[49030] = 0;
// bram[49031] = 0;
// bram[49032] = 5;
// bram[49033] = 15;
// bram[49034] = 29;
// bram[49035] = 46;
// bram[49036] = 67;
// bram[49037] = 89;
// bram[49038] = 113;
// bram[49039] = 138;
// bram[49040] = 162;
// bram[49041] = 185;
// bram[49042] = 205;
// bram[49043] = 223;
// bram[49044] = 237;
// bram[49045] = 247;
// bram[49046] = 252;
// bram[49047] = 253;
// bram[49048] = 249;
// bram[49049] = 241;
// bram[49050] = 228;
// bram[49051] = 211;
// bram[49052] = 191;
// bram[49053] = 169;
// bram[49054] = 145;
// bram[49055] = 121;
// bram[49056] = 96;
// bram[49057] = 73;
// bram[49058] = 52;
// bram[49059] = 34;
// bram[49060] = 19;
// bram[49061] = 8;
// bram[49062] = 1;
// bram[49063] = 0;
// bram[49064] = 2;
// bram[49065] = 10;
// bram[49066] = 22;
// bram[49067] = 38;
// bram[49068] = 57;
// bram[49069] = 79;
// bram[49070] = 102;
// bram[49071] = 127;
// bram[49072] = 151;
// bram[49073] = 175;
// bram[49074] = 196;
// bram[49075] = 215;
// bram[49076] = 231;
// bram[49077] = 243;
// bram[49078] = 251;
// bram[49079] = 253;
// bram[49080] = 252;
// bram[49081] = 245;
// bram[49082] = 234;
// bram[49083] = 219;
// bram[49084] = 201;
// bram[49085] = 179;
// bram[49086] = 156;
// bram[49087] = 132;
// bram[49088] = 107;
// bram[49089] = 84;
// bram[49090] = 61;
// bram[49091] = 42;
// bram[49092] = 25;
// bram[49093] = 12;
// bram[49094] = 4;
// bram[49095] = 0;
// bram[49096] = 1;
// bram[49097] = 6;
// bram[49098] = 16;
// bram[49099] = 30;
// bram[49100] = 48;
// bram[49101] = 69;
// bram[49102] = 91;
// bram[49103] = 115;
// bram[49104] = 140;
// bram[49105] = 164;
// bram[49106] = 187;
// bram[49107] = 207;
// bram[49108] = 224;
// bram[49109] = 238;
// bram[49110] = 248;
// bram[49111] = 253;
// bram[49112] = 253;
// bram[49113] = 249;
// bram[49114] = 240;
// bram[49115] = 226;
// bram[49116] = 209;
// bram[49117] = 189;
// bram[49118] = 167;
// bram[49119] = 143;
// bram[49120] = 119;
// bram[49121] = 94;
// bram[49122] = 71;
// bram[49123] = 50;
// bram[49124] = 32;
// bram[49125] = 18;
// bram[49126] = 7;
// bram[49127] = 1;
// bram[49128] = 0;
// bram[49129] = 3;
// bram[49130] = 11;
// bram[49131] = 23;
// bram[49132] = 39;
// bram[49133] = 59;
// bram[49134] = 81;
// bram[49135] = 104;
// bram[49136] = 129;
// bram[49137] = 153;
// bram[49138] = 177;
// bram[49139] = 198;
// bram[49140] = 217;
// bram[49141] = 232;
// bram[49142] = 244;
// bram[49143] = 251;
// bram[49144] = 253;
// bram[49145] = 251;
// bram[49146] = 244;
// bram[49147] = 233;
// bram[49148] = 218;
// bram[49149] = 199;
// bram[49150] = 177;
// bram[49151] = 154;
// bram[49152] = 130;
// bram[49153] = 105;
// bram[49154] = 82;
// bram[49155] = 60;
// bram[49156] = 40;
// bram[49157] = 24;
// bram[49158] = 11;
// bram[49159] = 3;
// bram[49160] = 0;
// bram[49161] = 1;
// bram[49162] = 7;
// bram[49163] = 17;
// bram[49164] = 32;
// bram[49165] = 50;
// bram[49166] = 71;
// bram[49167] = 94;
// bram[49168] = 118;
// bram[49169] = 142;
// bram[49170] = 166;
// bram[49171] = 189;
// bram[49172] = 209;
// bram[49173] = 226;
// bram[49174] = 239;
// bram[49175] = 248;
// bram[49176] = 253;
// bram[49177] = 253;
// bram[49178] = 248;
// bram[49179] = 239;
// bram[49180] = 225;
// bram[49181] = 208;
// bram[49182] = 187;
// bram[49183] = 165;
// bram[49184] = 141;
// bram[49185] = 116;
// bram[49186] = 92;
// bram[49187] = 69;
// bram[49188] = 49;
// bram[49189] = 31;
// bram[49190] = 16;
// bram[49191] = 6;
// bram[49192] = 1;
// bram[49193] = 0;
// bram[49194] = 4;
// bram[49195] = 12;
// bram[49196] = 25;
// bram[49197] = 41;
// bram[49198] = 61;
// bram[49199] = 83;
// bram[49200] = 107;
// bram[49201] = 131;
// bram[49202] = 155;
// bram[49203] = 179;
// bram[49204] = 200;
// bram[49205] = 219;
// bram[49206] = 234;
// bram[49207] = 245;
// bram[49208] = 251;
// bram[49209] = 253;
// bram[49210] = 251;
// bram[49211] = 243;
// bram[49212] = 232;
// bram[49213] = 216;
// bram[49214] = 197;
// bram[49215] = 175;
// bram[49216] = 152;
// bram[49217] = 127;
// bram[49218] = 103;
// bram[49219] = 79;
// bram[49220] = 58;
// bram[49221] = 38;
// bram[49222] = 22;
// bram[49223] = 10;
// bram[49224] = 3;
// bram[49225] = 0;
// bram[49226] = 1;
// bram[49227] = 8;
// bram[49228] = 18;
// bram[49229] = 33;
// bram[49230] = 51;
// bram[49231] = 73;
// bram[49232] = 96;
// bram[49233] = 120;
// bram[49234] = 144;
// bram[49235] = 168;
// bram[49236] = 191;
// bram[49237] = 211;
// bram[49238] = 227;
// bram[49239] = 240;
// bram[49240] = 249;
// bram[49241] = 253;
// bram[49242] = 253;
// bram[49243] = 247;
// bram[49244] = 238;
// bram[49245] = 224;
// bram[49246] = 206;
// bram[49247] = 185;
// bram[49248] = 163;
// bram[49249] = 139;
// bram[49250] = 114;
// bram[49251] = 90;
// bram[49252] = 67;
// bram[49253] = 47;
// bram[49254] = 29;
// bram[49255] = 15;
// bram[49256] = 6;
// bram[49257] = 0;
// bram[49258] = 0;
// bram[49259] = 4;
// bram[49260] = 13;
// bram[49261] = 26;
// bram[49262] = 43;
// bram[49263] = 63;
// bram[49264] = 85;
// bram[49265] = 109;
// bram[49266] = 133;
// bram[49267] = 158;
// bram[49268] = 181;
// bram[49269] = 202;
// bram[49270] = 220;
// bram[49271] = 235;
// bram[49272] = 246;
// bram[49273] = 252;
// bram[49274] = 253;
// bram[49275] = 250;
// bram[49276] = 242;
// bram[49277] = 230;
// bram[49278] = 214;
// bram[49279] = 195;
// bram[49280] = 173;
// bram[49281] = 150;
// bram[49282] = 125;
// bram[49283] = 101;
// bram[49284] = 77;
// bram[49285] = 56;
// bram[49286] = 37;
// bram[49287] = 21;
// bram[49288] = 9;
// bram[49289] = 2;
// bram[49290] = 0;
// bram[49291] = 2;
// bram[49292] = 8;
// bram[49293] = 20;
// bram[49294] = 35;
// bram[49295] = 53;
// bram[49296] = 75;
// bram[49297] = 98;
// bram[49298] = 122;
// bram[49299] = 147;
// bram[49300] = 170;
// bram[49301] = 193;
// bram[49302] = 212;
// bram[49303] = 229;
// bram[49304] = 241;
// bram[49305] = 250;
// bram[49306] = 253;
// bram[49307] = 252;
// bram[49308] = 247;
// bram[49309] = 236;
// bram[49310] = 222;
// bram[49311] = 204;
// bram[49312] = 183;
// bram[49313] = 161;
// bram[49314] = 136;
// bram[49315] = 112;
// bram[49316] = 88;
// bram[49317] = 65;
// bram[49318] = 45;
// bram[49319] = 28;
// bram[49320] = 14;
// bram[49321] = 5;
// bram[49322] = 0;
// bram[49323] = 0;
// bram[49324] = 5;
// bram[49325] = 14;
// bram[49326] = 27;
// bram[49327] = 44;
// bram[49328] = 65;
// bram[49329] = 87;
// bram[49330] = 111;
// bram[49331] = 136;
// bram[49332] = 160;
// bram[49333] = 183;
// bram[49334] = 204;
// bram[49335] = 222;
// bram[49336] = 236;
// bram[49337] = 246;
// bram[49338] = 252;
// bram[49339] = 253;
// bram[49340] = 250;
// bram[49341] = 242;
// bram[49342] = 229;
// bram[49343] = 213;
// bram[49344] = 193;
// bram[49345] = 171;
// bram[49346] = 147;
// bram[49347] = 123;
// bram[49348] = 99;
// bram[49349] = 75;
// bram[49350] = 54;
// bram[49351] = 35;
// bram[49352] = 20;
// bram[49353] = 9;
// bram[49354] = 2;
// bram[49355] = 0;
// bram[49356] = 2;
// bram[49357] = 9;
// bram[49358] = 21;
// bram[49359] = 36;
// bram[49360] = 55;
// bram[49361] = 77;
// bram[49362] = 100;
// bram[49363] = 124;
// bram[49364] = 149;
// bram[49365] = 173;
// bram[49366] = 194;
// bram[49367] = 214;
// bram[49368] = 230;
// bram[49369] = 242;
// bram[49370] = 250;
// bram[49371] = 253;
// bram[49372] = 252;
// bram[49373] = 246;
// bram[49374] = 235;
// bram[49375] = 221;
// bram[49376] = 202;
// bram[49377] = 181;
// bram[49378] = 158;
// bram[49379] = 134;
// bram[49380] = 110;
// bram[49381] = 86;
// bram[49382] = 63;
// bram[49383] = 43;
// bram[49384] = 26;
// bram[49385] = 13;
// bram[49386] = 4;
// bram[49387] = 0;
// bram[49388] = 0;
// bram[49389] = 5;
// bram[49390] = 15;
// bram[49391] = 29;
// bram[49392] = 46;
// bram[49393] = 67;
// bram[49394] = 89;
// bram[49395] = 113;
// bram[49396] = 138;
// bram[49397] = 162;
// bram[49398] = 185;
// bram[49399] = 205;
// bram[49400] = 223;
// bram[49401] = 237;
// bram[49402] = 247;
// bram[49403] = 252;
// bram[49404] = 253;
// bram[49405] = 249;
// bram[49406] = 241;
// bram[49407] = 228;
// bram[49408] = 211;
// bram[49409] = 191;
// bram[49410] = 169;
// bram[49411] = 145;
// bram[49412] = 121;
// bram[49413] = 96;
// bram[49414] = 73;
// bram[49415] = 52;
// bram[49416] = 34;
// bram[49417] = 19;
// bram[49418] = 8;
// bram[49419] = 1;
// bram[49420] = 0;
// bram[49421] = 2;
// bram[49422] = 10;
// bram[49423] = 22;
// bram[49424] = 38;
// bram[49425] = 57;
// bram[49426] = 79;
// bram[49427] = 102;
// bram[49428] = 127;
// bram[49429] = 151;
// bram[49430] = 175;
// bram[49431] = 196;
// bram[49432] = 215;
// bram[49433] = 231;
// bram[49434] = 243;
// bram[49435] = 251;
// bram[49436] = 253;
// bram[49437] = 252;
// bram[49438] = 245;
// bram[49439] = 234;
// bram[49440] = 219;
// bram[49441] = 201;
// bram[49442] = 179;
// bram[49443] = 156;
// bram[49444] = 132;
// bram[49445] = 107;
// bram[49446] = 84;
// bram[49447] = 61;
// bram[49448] = 42;
// bram[49449] = 25;
// bram[49450] = 12;
// bram[49451] = 4;
// bram[49452] = 0;
// bram[49453] = 1;
// bram[49454] = 6;
// bram[49455] = 16;
// bram[49456] = 30;
// bram[49457] = 48;
// bram[49458] = 69;
// bram[49459] = 91;
// bram[49460] = 116;
// bram[49461] = 140;
// bram[49462] = 164;
// bram[49463] = 187;
// bram[49464] = 207;
// bram[49465] = 225;
// bram[49466] = 238;
// bram[49467] = 248;
// bram[49468] = 253;
// bram[49469] = 253;
// bram[49470] = 249;
// bram[49471] = 240;
// bram[49472] = 226;
// bram[49473] = 209;
// bram[49474] = 189;
// bram[49475] = 167;
// bram[49476] = 143;
// bram[49477] = 118;
// bram[49478] = 94;
// bram[49479] = 71;
// bram[49480] = 50;
// bram[49481] = 32;
// bram[49482] = 18;
// bram[49483] = 7;
// bram[49484] = 1;
// bram[49485] = 0;
// bram[49486] = 3;
// bram[49487] = 11;
// bram[49488] = 23;
// bram[49489] = 39;
// bram[49490] = 59;
// bram[49491] = 81;
// bram[49492] = 104;
// bram[49493] = 129;
// bram[49494] = 153;
// bram[49495] = 177;
// bram[49496] = 198;
// bram[49497] = 217;
// bram[49498] = 232;
// bram[49499] = 244;
// bram[49500] = 251;
// bram[49501] = 253;
// bram[49502] = 251;
// bram[49503] = 244;
// bram[49504] = 233;
// bram[49505] = 218;
// bram[49506] = 199;
// bram[49507] = 177;
// bram[49508] = 154;
// bram[49509] = 130;
// bram[49510] = 105;
// bram[49511] = 81;
// bram[49512] = 59;
// bram[49513] = 40;
// bram[49514] = 24;
// bram[49515] = 11;
// bram[49516] = 3;
// bram[49517] = 0;
// bram[49518] = 1;
// bram[49519] = 7;
// bram[49520] = 17;
// bram[49521] = 32;
// bram[49522] = 50;
// bram[49523] = 71;
// bram[49524] = 94;
// bram[49525] = 118;
// bram[49526] = 142;
// bram[49527] = 166;
// bram[49528] = 189;
// bram[49529] = 209;
// bram[49530] = 226;
// bram[49531] = 239;
// bram[49532] = 248;
// bram[49533] = 253;
// bram[49534] = 253;
// bram[49535] = 248;
// bram[49536] = 239;
// bram[49537] = 225;
// bram[49538] = 208;
// bram[49539] = 187;
// bram[49540] = 165;
// bram[49541] = 141;
// bram[49542] = 116;
// bram[49543] = 92;
// bram[49544] = 69;
// bram[49545] = 48;
// bram[49546] = 31;
// bram[49547] = 16;
// bram[49548] = 6;
// bram[49549] = 1;
// bram[49550] = 0;
// bram[49551] = 4;
// bram[49552] = 12;
// bram[49553] = 25;
// bram[49554] = 41;
// bram[49555] = 61;
// bram[49556] = 83;
// bram[49557] = 107;
// bram[49558] = 131;
// bram[49559] = 156;
// bram[49560] = 179;
// bram[49561] = 200;
// bram[49562] = 219;
// bram[49563] = 234;
// bram[49564] = 245;
// bram[49565] = 251;
// bram[49566] = 253;
// bram[49567] = 251;
// bram[49568] = 243;
// bram[49569] = 232;
// bram[49570] = 216;
// bram[49571] = 197;
// bram[49572] = 175;
// bram[49573] = 152;
// bram[49574] = 127;
// bram[49575] = 103;
// bram[49576] = 79;
// bram[49577] = 58;
// bram[49578] = 38;
// bram[49579] = 22;
// bram[49580] = 10;
// bram[49581] = 3;
// bram[49582] = 0;
// bram[49583] = 1;
// bram[49584] = 8;
// bram[49585] = 18;
// bram[49586] = 33;
// bram[49587] = 51;
// bram[49588] = 73;
// bram[49589] = 96;
// bram[49590] = 120;
// bram[49591] = 145;
// bram[49592] = 168;
// bram[49593] = 191;
// bram[49594] = 211;
// bram[49595] = 227;
// bram[49596] = 240;
// bram[49597] = 249;
// bram[49598] = 253;
// bram[49599] = 253;
// bram[49600] = 247;
// bram[49601] = 237;
// bram[49602] = 224;
// bram[49603] = 206;
// bram[49604] = 185;
// bram[49605] = 163;
// bram[49606] = 139;
// bram[49607] = 114;
// bram[49608] = 90;
// bram[49609] = 67;
// bram[49610] = 47;
// bram[49611] = 29;
// bram[49612] = 15;
// bram[49613] = 6;
// bram[49614] = 0;
// bram[49615] = 0;
// bram[49616] = 4;
// bram[49617] = 13;
// bram[49618] = 26;
// bram[49619] = 43;
// bram[49620] = 63;
// bram[49621] = 85;
// bram[49622] = 109;
// bram[49623] = 133;
// bram[49624] = 158;
// bram[49625] = 181;
// bram[49626] = 202;
// bram[49627] = 220;
// bram[49628] = 235;
// bram[49629] = 246;
// bram[49630] = 252;
// bram[49631] = 253;
// bram[49632] = 250;
// bram[49633] = 242;
// bram[49634] = 230;
// bram[49635] = 214;
// bram[49636] = 195;
// bram[49637] = 173;
// bram[49638] = 150;
// bram[49639] = 125;
// bram[49640] = 101;
// bram[49641] = 77;
// bram[49642] = 56;
// bram[49643] = 37;
// bram[49644] = 21;
// bram[49645] = 9;
// bram[49646] = 2;
// bram[49647] = 0;
// bram[49648] = 2;
// bram[49649] = 8;
// bram[49650] = 20;
// bram[49651] = 35;
// bram[49652] = 53;
// bram[49653] = 75;
// bram[49654] = 98;
// bram[49655] = 122;
// bram[49656] = 147;
// bram[49657] = 171;
// bram[49658] = 193;
// bram[49659] = 212;
// bram[49660] = 229;
// bram[49661] = 241;
// bram[49662] = 250;
// bram[49663] = 253;
// bram[49664] = 252;
// bram[49665] = 247;
// bram[49666] = 236;
// bram[49667] = 222;
// bram[49668] = 204;
// bram[49669] = 183;
// bram[49670] = 160;
// bram[49671] = 136;
// bram[49672] = 112;
// bram[49673] = 88;
// bram[49674] = 65;
// bram[49675] = 45;
// bram[49676] = 28;
// bram[49677] = 14;
// bram[49678] = 5;
// bram[49679] = 0;
// bram[49680] = 0;
// bram[49681] = 5;
// bram[49682] = 14;
// bram[49683] = 27;
// bram[49684] = 44;
// bram[49685] = 65;
// bram[49686] = 87;
// bram[49687] = 111;
// bram[49688] = 136;
// bram[49689] = 160;
// bram[49690] = 183;
// bram[49691] = 204;
// bram[49692] = 222;
// bram[49693] = 236;
// bram[49694] = 246;
// bram[49695] = 252;
// bram[49696] = 253;
// bram[49697] = 250;
// bram[49698] = 242;
// bram[49699] = 229;
// bram[49700] = 213;
// bram[49701] = 193;
// bram[49702] = 171;
// bram[49703] = 147;
// bram[49704] = 123;
// bram[49705] = 99;
// bram[49706] = 75;
// bram[49707] = 54;
// bram[49708] = 35;
// bram[49709] = 20;
// bram[49710] = 9;
// bram[49711] = 2;
// bram[49712] = 0;
// bram[49713] = 2;
// bram[49714] = 9;
// bram[49715] = 21;
// bram[49716] = 36;
// bram[49717] = 55;
// bram[49718] = 77;
// bram[49719] = 100;
// bram[49720] = 125;
// bram[49721] = 149;
// bram[49722] = 173;
// bram[49723] = 195;
// bram[49724] = 214;
// bram[49725] = 230;
// bram[49726] = 242;
// bram[49727] = 250;
// bram[49728] = 253;
// bram[49729] = 252;
// bram[49730] = 246;
// bram[49731] = 235;
// bram[49732] = 221;
// bram[49733] = 202;
// bram[49734] = 181;
// bram[49735] = 158;
// bram[49736] = 134;
// bram[49737] = 110;
// bram[49738] = 86;
// bram[49739] = 63;
// bram[49740] = 43;
// bram[49741] = 26;
// bram[49742] = 13;
// bram[49743] = 4;
// bram[49744] = 0;
// bram[49745] = 0;
// bram[49746] = 5;
// bram[49747] = 15;
// bram[49748] = 29;
// bram[49749] = 46;
// bram[49750] = 67;
// bram[49751] = 89;
// bram[49752] = 113;
// bram[49753] = 138;
// bram[49754] = 162;
// bram[49755] = 185;
// bram[49756] = 205;
// bram[49757] = 223;
// bram[49758] = 237;
// bram[49759] = 247;
// bram[49760] = 252;
// bram[49761] = 253;
// bram[49762] = 249;
// bram[49763] = 241;
// bram[49764] = 228;
// bram[49765] = 211;
// bram[49766] = 191;
// bram[49767] = 169;
// bram[49768] = 145;
// bram[49769] = 121;
// bram[49770] = 96;
// bram[49771] = 73;
// bram[49772] = 52;
// bram[49773] = 34;
// bram[49774] = 19;
// bram[49775] = 8;
// bram[49776] = 1;
// bram[49777] = 0;
// bram[49778] = 2;
// bram[49779] = 10;
// bram[49780] = 22;
// bram[49781] = 38;
// bram[49782] = 57;
// bram[49783] = 79;
// bram[49784] = 102;
// bram[49785] = 127;
// bram[49786] = 151;
// bram[49787] = 175;
// bram[49788] = 196;
// bram[49789] = 215;
// bram[49790] = 231;
// bram[49791] = 243;
// bram[49792] = 251;
// bram[49793] = 253;
// bram[49794] = 252;
// bram[49795] = 245;
// bram[49796] = 234;
// bram[49797] = 219;
// bram[49798] = 201;
// bram[49799] = 179;
// bram[49800] = 156;
// bram[49801] = 132;
// bram[49802] = 107;
// bram[49803] = 84;
// bram[49804] = 61;
// bram[49805] = 42;
// bram[49806] = 25;
// bram[49807] = 12;
// bram[49808] = 4;
// bram[49809] = 0;
// bram[49810] = 1;
// bram[49811] = 6;
// bram[49812] = 16;
// bram[49813] = 30;
// bram[49814] = 48;
// bram[49815] = 69;
// bram[49816] = 91;
// bram[49817] = 116;
// bram[49818] = 140;
// bram[49819] = 164;
// bram[49820] = 187;
// bram[49821] = 207;
// bram[49822] = 225;
// bram[49823] = 238;
// bram[49824] = 248;
// bram[49825] = 253;
// bram[49826] = 253;
// bram[49827] = 249;
// bram[49828] = 240;
// bram[49829] = 226;
// bram[49830] = 209;
// bram[49831] = 189;
// bram[49832] = 167;
// bram[49833] = 143;
// bram[49834] = 118;
// bram[49835] = 94;
// bram[49836] = 71;
// bram[49837] = 50;
// bram[49838] = 32;
// bram[49839] = 18;
// bram[49840] = 7;
// bram[49841] = 1;
// bram[49842] = 0;
// bram[49843] = 3;
// bram[49844] = 11;
// bram[49845] = 23;
// bram[49846] = 39;
// bram[49847] = 59;
// bram[49848] = 81;
// bram[49849] = 105;
// bram[49850] = 129;
// bram[49851] = 153;
// bram[49852] = 177;
// bram[49853] = 198;
// bram[49854] = 217;
// bram[49855] = 233;
// bram[49856] = 244;
// bram[49857] = 251;
// bram[49858] = 253;
// bram[49859] = 251;
// bram[49860] = 244;
// bram[49861] = 233;
// bram[49862] = 217;
// bram[49863] = 199;
// bram[49864] = 177;
// bram[49865] = 154;
// bram[49866] = 130;
// bram[49867] = 105;
// bram[49868] = 81;
// bram[49869] = 59;
// bram[49870] = 40;
// bram[49871] = 24;
// bram[49872] = 11;
// bram[49873] = 3;
// bram[49874] = 0;
// bram[49875] = 1;
// bram[49876] = 7;
// bram[49877] = 17;
// bram[49878] = 32;
// bram[49879] = 50;
// bram[49880] = 71;
// bram[49881] = 94;
// bram[49882] = 118;
// bram[49883] = 142;
// bram[49884] = 166;
// bram[49885] = 189;
// bram[49886] = 209;
// bram[49887] = 226;
// bram[49888] = 239;
// bram[49889] = 248;
// bram[49890] = 253;
// bram[49891] = 253;
// bram[49892] = 248;
// bram[49893] = 239;
// bram[49894] = 225;
// bram[49895] = 208;
// bram[49896] = 187;
// bram[49897] = 165;
// bram[49898] = 141;
// bram[49899] = 116;
// bram[49900] = 92;
// bram[49901] = 69;
// bram[49902] = 48;
// bram[49903] = 31;
// bram[49904] = 16;
// bram[49905] = 6;
// bram[49906] = 1;
// bram[49907] = 0;
// bram[49908] = 4;
// bram[49909] = 12;
// bram[49910] = 25;
// bram[49911] = 41;
// bram[49912] = 61;
// bram[49913] = 83;
// bram[49914] = 107;
// bram[49915] = 131;
// bram[49916] = 156;
// bram[49917] = 179;
// bram[49918] = 200;
// bram[49919] = 219;
// bram[49920] = 234;
// bram[49921] = 245;
// bram[49922] = 251;
// bram[49923] = 253;
// bram[49924] = 251;
// bram[49925] = 243;
// bram[49926] = 232;
// bram[49927] = 216;
// bram[49928] = 197;
// bram[49929] = 175;
// bram[49930] = 152;
// bram[49931] = 127;
// bram[49932] = 103;
// bram[49933] = 79;
// bram[49934] = 58;
// bram[49935] = 38;
// bram[49936] = 22;
// bram[49937] = 10;
// bram[49938] = 3;
// bram[49939] = 0;
// bram[49940] = 1;
// bram[49941] = 8;
// bram[49942] = 18;
// bram[49943] = 33;
// bram[49944] = 52;
// bram[49945] = 73;
// bram[49946] = 96;
// bram[49947] = 120;
// bram[49948] = 145;
// bram[49949] = 168;
// bram[49950] = 191;
// bram[49951] = 211;
// bram[49952] = 227;
// bram[49953] = 240;
// bram[49954] = 249;
// bram[49955] = 253;
// bram[49956] = 253;
// bram[49957] = 247;
// bram[49958] = 237;
// bram[49959] = 223;
// bram[49960] = 206;
// bram[49961] = 185;
// bram[49962] = 163;
// bram[49963] = 139;
// bram[49964] = 114;
// bram[49965] = 90;
// bram[49966] = 67;
// bram[49967] = 47;
// bram[49968] = 29;
// bram[49969] = 15;
// bram[49970] = 6;
// bram[49971] = 0;
// bram[49972] = 0;
// bram[49973] = 4;
// bram[49974] = 13;
// bram[49975] = 26;
// bram[49976] = 43;
// bram[49977] = 63;
// bram[49978] = 85;
// bram[49979] = 109;
// bram[49980] = 133;
// bram[49981] = 158;
// bram[49982] = 181;
// bram[49983] = 202;
// bram[49984] = 220;
// bram[49985] = 235;
// bram[49986] = 246;
// bram[49987] = 252;
// bram[49988] = 253;
// bram[49989] = 250;
// bram[49990] = 242;
// bram[49991] = 230;
// bram[49992] = 214;
// bram[49993] = 195;
// bram[49994] = 173;
// bram[49995] = 150;
// bram[49996] = 125;
// bram[49997] = 101;
// bram[49998] = 77;
// bram[49999] = 56;
// bram[50000] = 37;
// bram[50001] = 21;
// bram[50002] = 9;
// bram[50003] = 2;
// bram[50004] = 0;
// bram[50005] = 2;
// bram[50006] = 8;
// bram[50007] = 20;
// bram[50008] = 35;
// bram[50009] = 53;
// bram[50010] = 75;
// bram[50011] = 98;
// bram[50012] = 122;
// bram[50013] = 147;
// bram[50014] = 171;
// bram[50015] = 193;
// bram[50016] = 212;
// bram[50017] = 229;
// bram[50018] = 241;
// bram[50019] = 250;
// bram[50020] = 253;
// bram[50021] = 252;
// bram[50022] = 247;
// bram[50023] = 236;
// bram[50024] = 222;
// bram[50025] = 204;
// bram[50026] = 183;
// bram[50027] = 160;
// bram[50028] = 136;
// bram[50029] = 112;
// bram[50030] = 88;
// bram[50031] = 65;
// bram[50032] = 45;
// bram[50033] = 28;
// bram[50034] = 14;
// bram[50035] = 5;
// bram[50036] = 0;
// bram[50037] = 0;
// bram[50038] = 5;
// bram[50039] = 14;
// bram[50040] = 27;
// bram[50041] = 45;
// bram[50042] = 65;
// bram[50043] = 87;
// bram[50044] = 111;
// bram[50045] = 136;
// bram[50046] = 160;
// bram[50047] = 183;
// bram[50048] = 204;
// bram[50049] = 222;
// bram[50050] = 236;
// bram[50051] = 246;
// bram[50052] = 252;
// bram[50053] = 253;
// bram[50054] = 250;
// bram[50055] = 242;
// bram[50056] = 229;
// bram[50057] = 213;
// bram[50058] = 193;
// bram[50059] = 171;
// bram[50060] = 147;
// bram[50061] = 123;
// bram[50062] = 99;
// bram[50063] = 75;
// bram[50064] = 54;
// bram[50065] = 35;
// bram[50066] = 20;
// bram[50067] = 9;
// bram[50068] = 2;
// bram[50069] = 0;
// bram[50070] = 2;
// bram[50071] = 9;
// bram[50072] = 21;
// bram[50073] = 36;
// bram[50074] = 55;
// bram[50075] = 77;
// bram[50076] = 100;
// bram[50077] = 125;
// bram[50078] = 149;
// bram[50079] = 173;
// bram[50080] = 195;
// bram[50081] = 214;
// bram[50082] = 230;
// bram[50083] = 242;
// bram[50084] = 250;
// bram[50085] = 253;
// bram[50086] = 252;
// bram[50087] = 246;
// bram[50088] = 235;
// bram[50089] = 221;
// bram[50090] = 202;
// bram[50091] = 181;
// bram[50092] = 158;
// bram[50093] = 134;
// bram[50094] = 109;
// bram[50095] = 86;
// bram[50096] = 63;
// bram[50097] = 43;
// bram[50098] = 26;
// bram[50099] = 13;
// bram[50100] = 4;
// bram[50101] = 0;
// bram[50102] = 0;
// bram[50103] = 5;
// bram[50104] = 15;
// bram[50105] = 29;
// bram[50106] = 46;
// bram[50107] = 67;
// bram[50108] = 89;
// bram[50109] = 113;
// bram[50110] = 138;
// bram[50111] = 162;
// bram[50112] = 185;
// bram[50113] = 205;
// bram[50114] = 223;
// bram[50115] = 237;
// bram[50116] = 247;
// bram[50117] = 253;
// bram[50118] = 253;
// bram[50119] = 249;
// bram[50120] = 241;
// bram[50121] = 228;
// bram[50122] = 211;
// bram[50123] = 191;
// bram[50124] = 169;
// bram[50125] = 145;
// bram[50126] = 121;
// bram[50127] = 96;
// bram[50128] = 73;
// bram[50129] = 52;
// bram[50130] = 34;
// bram[50131] = 19;
// bram[50132] = 8;
// bram[50133] = 1;
// bram[50134] = 0;
// bram[50135] = 3;
// bram[50136] = 10;
// bram[50137] = 22;
// bram[50138] = 38;
// bram[50139] = 57;
// bram[50140] = 79;
// bram[50141] = 102;
// bram[50142] = 127;
// bram[50143] = 151;
// bram[50144] = 175;
// bram[50145] = 196;
// bram[50146] = 216;
// bram[50147] = 231;
// bram[50148] = 243;
// bram[50149] = 251;
// bram[50150] = 253;
// bram[50151] = 252;
// bram[50152] = 245;
// bram[50153] = 234;
// bram[50154] = 219;
// bram[50155] = 201;
// bram[50156] = 179;
// bram[50157] = 156;
// bram[50158] = 132;
// bram[50159] = 107;
// bram[50160] = 83;
// bram[50161] = 61;
// bram[50162] = 42;
// bram[50163] = 25;
// bram[50164] = 12;
// bram[50165] = 4;
// bram[50166] = 0;
// bram[50167] = 1;
// bram[50168] = 6;
// bram[50169] = 16;
// bram[50170] = 30;
// bram[50171] = 48;
// bram[50172] = 69;
// bram[50173] = 91;
// bram[50174] = 116;
// bram[50175] = 140;
// bram[50176] = 164;
// bram[50177] = 187;
// bram[50178] = 207;
// bram[50179] = 225;
// bram[50180] = 238;
// bram[50181] = 248;
// bram[50182] = 253;
// bram[50183] = 253;
// bram[50184] = 249;
// bram[50185] = 240;
// bram[50186] = 226;
// bram[50187] = 209;
// bram[50188] = 189;
// bram[50189] = 167;
// bram[50190] = 143;
// bram[50191] = 118;
// bram[50192] = 94;
// bram[50193] = 71;
// bram[50194] = 50;
// bram[50195] = 32;
// bram[50196] = 17;
// bram[50197] = 7;
// bram[50198] = 1;
// bram[50199] = 0;
// bram[50200] = 3;
// bram[50201] = 11;
// bram[50202] = 23;
// bram[50203] = 40;
// bram[50204] = 59;
// bram[50205] = 81;
// bram[50206] = 105;
// bram[50207] = 129;
// bram[50208] = 153;
// bram[50209] = 177;
// bram[50210] = 198;
// bram[50211] = 217;
// bram[50212] = 233;
// bram[50213] = 244;
// bram[50214] = 251;
// bram[50215] = 253;
// bram[50216] = 251;
// bram[50217] = 244;
// bram[50218] = 233;
// bram[50219] = 217;
// bram[50220] = 199;
// bram[50221] = 177;
// bram[50222] = 154;
// bram[50223] = 130;
// bram[50224] = 105;
// bram[50225] = 81;
// bram[50226] = 59;
// bram[50227] = 40;
// bram[50228] = 24;
// bram[50229] = 11;
// bram[50230] = 3;
// bram[50231] = 0;
// bram[50232] = 1;
// bram[50233] = 7;
// bram[50234] = 17;
// bram[50235] = 32;
// bram[50236] = 50;
// bram[50237] = 71;
// bram[50238] = 94;
// bram[50239] = 118;
// bram[50240] = 142;
// bram[50241] = 166;
// bram[50242] = 189;
// bram[50243] = 209;
// bram[50244] = 226;
// bram[50245] = 239;
// bram[50246] = 248;
// bram[50247] = 253;
// bram[50248] = 253;
// bram[50249] = 248;
// bram[50250] = 239;
// bram[50251] = 225;
// bram[50252] = 208;
// bram[50253] = 187;
// bram[50254] = 165;
// bram[50255] = 141;
// bram[50256] = 116;
// bram[50257] = 92;
// bram[50258] = 69;
// bram[50259] = 48;
// bram[50260] = 31;
// bram[50261] = 16;
// bram[50262] = 6;
// bram[50263] = 1;
// bram[50264] = 0;
// bram[50265] = 4;
// bram[50266] = 12;
// bram[50267] = 25;
// bram[50268] = 41;
// bram[50269] = 61;
// bram[50270] = 83;
// bram[50271] = 107;
// bram[50272] = 131;
// bram[50273] = 156;
// bram[50274] = 179;
// bram[50275] = 200;
// bram[50276] = 219;
// bram[50277] = 234;
// bram[50278] = 245;
// bram[50279] = 251;
// bram[50280] = 253;
// bram[50281] = 251;
// bram[50282] = 243;
// bram[50283] = 232;
// bram[50284] = 216;
// bram[50285] = 197;
// bram[50286] = 175;
// bram[50287] = 152;
// bram[50288] = 127;
// bram[50289] = 103;
// bram[50290] = 79;
// bram[50291] = 57;
// bram[50292] = 38;
// bram[50293] = 22;
// bram[50294] = 10;
// bram[50295] = 3;
// bram[50296] = 0;
// bram[50297] = 1;
// bram[50298] = 8;
// bram[50299] = 18;
// bram[50300] = 33;
// bram[50301] = 52;
// bram[50302] = 73;
// bram[50303] = 96;
// bram[50304] = 120;
// bram[50305] = 145;
// bram[50306] = 168;
// bram[50307] = 191;
// bram[50308] = 211;
// bram[50309] = 227;
// bram[50310] = 240;
// bram[50311] = 249;
// bram[50312] = 253;
// bram[50313] = 253;
// bram[50314] = 247;
// bram[50315] = 237;
// bram[50316] = 223;
// bram[50317] = 206;
// bram[50318] = 185;
// bram[50319] = 163;
// bram[50320] = 138;
// bram[50321] = 114;
// bram[50322] = 90;
// bram[50323] = 67;
// bram[50324] = 47;
// bram[50325] = 29;
// bram[50326] = 15;
// bram[50327] = 6;
// bram[50328] = 0;
// bram[50329] = 0;
// bram[50330] = 4;
// bram[50331] = 13;
// bram[50332] = 26;
// bram[50333] = 43;
// bram[50334] = 63;
// bram[50335] = 85;
// bram[50336] = 109;
// bram[50337] = 134;
// bram[50338] = 158;
// bram[50339] = 181;
// bram[50340] = 202;
// bram[50341] = 220;
// bram[50342] = 235;
// bram[50343] = 246;
// bram[50344] = 252;
// bram[50345] = 253;
// bram[50346] = 250;
// bram[50347] = 242;
// bram[50348] = 230;
// bram[50349] = 214;
// bram[50350] = 195;
// bram[50351] = 173;
// bram[50352] = 150;
// bram[50353] = 125;
// bram[50354] = 101;
// bram[50355] = 77;
// bram[50356] = 56;
// bram[50357] = 37;
// bram[50358] = 21;
// bram[50359] = 9;
// bram[50360] = 2;
// bram[50361] = 0;
// bram[50362] = 2;
// bram[50363] = 8;
// bram[50364] = 20;
// bram[50365] = 35;
// bram[50366] = 53;
// bram[50367] = 75;
// bram[50368] = 98;
// bram[50369] = 122;
// bram[50370] = 147;
// bram[50371] = 171;
// bram[50372] = 193;
// bram[50373] = 212;
// bram[50374] = 229;
// bram[50375] = 241;
// bram[50376] = 250;
// bram[50377] = 253;
// bram[50378] = 252;
// bram[50379] = 247;
// bram[50380] = 236;
// bram[50381] = 222;
// bram[50382] = 204;
// bram[50383] = 183;
// bram[50384] = 160;
// bram[50385] = 136;
// bram[50386] = 112;
// bram[50387] = 88;
// bram[50388] = 65;
// bram[50389] = 45;
// bram[50390] = 28;
// bram[50391] = 14;
// bram[50392] = 5;
// bram[50393] = 0;
// bram[50394] = 0;
// bram[50395] = 5;
// bram[50396] = 14;
// bram[50397] = 27;
// bram[50398] = 45;
// bram[50399] = 65;
// bram[50400] = 87;
// bram[50401] = 111;
// bram[50402] = 136;
// bram[50403] = 160;
// bram[50404] = 183;
// bram[50405] = 204;
// bram[50406] = 222;
// bram[50407] = 236;
// bram[50408] = 246;
// bram[50409] = 252;
// bram[50410] = 253;
// bram[50411] = 250;
// bram[50412] = 241;
// bram[50413] = 229;
// bram[50414] = 213;
// bram[50415] = 193;
// bram[50416] = 171;
// bram[50417] = 147;
// bram[50418] = 123;
// bram[50419] = 98;
// bram[50420] = 75;
// bram[50421] = 54;
// bram[50422] = 35;
// bram[50423] = 20;
// bram[50424] = 9;
// bram[50425] = 2;
// bram[50426] = 0;
// bram[50427] = 2;
// bram[50428] = 9;
// bram[50429] = 21;
// bram[50430] = 36;
// bram[50431] = 55;
// bram[50432] = 77;
// bram[50433] = 100;
// bram[50434] = 125;
// bram[50435] = 149;
// bram[50436] = 173;
// bram[50437] = 195;
// bram[50438] = 214;
// bram[50439] = 230;
// bram[50440] = 242;
// bram[50441] = 250;
// bram[50442] = 253;
// bram[50443] = 252;
// bram[50444] = 246;
// bram[50445] = 235;
// bram[50446] = 221;
// bram[50447] = 202;
// bram[50448] = 181;
// bram[50449] = 158;
// bram[50450] = 134;
// bram[50451] = 109;
// bram[50452] = 86;
// bram[50453] = 63;
// bram[50454] = 43;
// bram[50455] = 26;
// bram[50456] = 13;
// bram[50457] = 4;
// bram[50458] = 0;
// bram[50459] = 0;
// bram[50460] = 5;
// bram[50461] = 15;
// bram[50462] = 29;
// bram[50463] = 46;
// bram[50464] = 67;
// bram[50465] = 89;
// bram[50466] = 113;
// bram[50467] = 138;
// bram[50468] = 162;
// bram[50469] = 185;
// bram[50470] = 206;
// bram[50471] = 223;
// bram[50472] = 237;
// bram[50473] = 247;
// bram[50474] = 253;
// bram[50475] = 253;
// bram[50476] = 249;
// bram[50477] = 241;
// bram[50478] = 228;
// bram[50479] = 211;
// bram[50480] = 191;
// bram[50481] = 169;
// bram[50482] = 145;
// bram[50483] = 121;
// bram[50484] = 96;
// bram[50485] = 73;
// bram[50486] = 52;
// bram[50487] = 34;
// bram[50488] = 19;
// bram[50489] = 8;
// bram[50490] = 1;
// bram[50491] = 0;
// bram[50492] = 3;
// bram[50493] = 10;
// bram[50494] = 22;
// bram[50495] = 38;
// bram[50496] = 57;
// bram[50497] = 79;
// bram[50498] = 102;
// bram[50499] = 127;
// bram[50500] = 151;
// bram[50501] = 175;
// bram[50502] = 196;
// bram[50503] = 216;
// bram[50504] = 231;
// bram[50505] = 243;
// bram[50506] = 251;
// bram[50507] = 253;
// bram[50508] = 252;
// bram[50509] = 245;
// bram[50510] = 234;
// bram[50511] = 219;
// bram[50512] = 201;
// bram[50513] = 179;
// bram[50514] = 156;
// bram[50515] = 132;
// bram[50516] = 107;
// bram[50517] = 83;
// bram[50518] = 61;
// bram[50519] = 42;
// bram[50520] = 25;
// bram[50521] = 12;
// bram[50522] = 4;
// bram[50523] = 0;
// bram[50524] = 1;
// bram[50525] = 6;
// bram[50526] = 16;
// bram[50527] = 30;
// bram[50528] = 48;
// bram[50529] = 69;
// bram[50530] = 92;
// bram[50531] = 116;
// bram[50532] = 140;
// bram[50533] = 164;
// bram[50534] = 187;
// bram[50535] = 207;
// bram[50536] = 225;
// bram[50537] = 238;
// bram[50538] = 248;
// bram[50539] = 253;
// bram[50540] = 253;
// bram[50541] = 249;
// bram[50542] = 240;
// bram[50543] = 226;
// bram[50544] = 209;
// bram[50545] = 189;
// bram[50546] = 167;
// bram[50547] = 143;
// bram[50548] = 118;
// bram[50549] = 94;
// bram[50550] = 71;
// bram[50551] = 50;
// bram[50552] = 32;
// bram[50553] = 17;
// bram[50554] = 7;
// bram[50555] = 1;
// bram[50556] = 0;
// bram[50557] = 3;
// bram[50558] = 11;
// bram[50559] = 23;
// bram[50560] = 40;
// bram[50561] = 59;
// bram[50562] = 81;
// bram[50563] = 105;
// bram[50564] = 129;
// bram[50565] = 153;
// bram[50566] = 177;
// bram[50567] = 198;
// bram[50568] = 217;
// bram[50569] = 233;
// bram[50570] = 244;
// bram[50571] = 251;
// bram[50572] = 253;
// bram[50573] = 251;
// bram[50574] = 244;
// bram[50575] = 233;
// bram[50576] = 217;
// bram[50577] = 199;
// bram[50578] = 177;
// bram[50579] = 154;
// bram[50580] = 129;
// bram[50581] = 105;
// bram[50582] = 81;
// bram[50583] = 59;
// bram[50584] = 40;
// bram[50585] = 24;
// bram[50586] = 11;
// bram[50587] = 3;
// bram[50588] = 0;
// bram[50589] = 1;
// bram[50590] = 7;
// bram[50591] = 17;
// bram[50592] = 32;
// bram[50593] = 50;
// bram[50594] = 71;
// bram[50595] = 94;
// bram[50596] = 118;
// bram[50597] = 142;
// bram[50598] = 166;
// bram[50599] = 189;
// bram[50600] = 209;
// bram[50601] = 226;
// bram[50602] = 239;
// bram[50603] = 248;
// bram[50604] = 253;
// bram[50605] = 253;
// bram[50606] = 248;
// bram[50607] = 238;
// bram[50608] = 225;
// bram[50609] = 208;
// bram[50610] = 187;
// bram[50611] = 165;
// bram[50612] = 141;
// bram[50613] = 116;
// bram[50614] = 92;
// bram[50615] = 69;
// bram[50616] = 48;
// bram[50617] = 31;
// bram[50618] = 16;
// bram[50619] = 6;
// bram[50620] = 1;
// bram[50621] = 0;
// bram[50622] = 4;
// bram[50623] = 12;
// bram[50624] = 25;
// bram[50625] = 41;
// bram[50626] = 61;
// bram[50627] = 83;
// bram[50628] = 107;
// bram[50629] = 131;
// bram[50630] = 156;
// bram[50631] = 179;
// bram[50632] = 200;
// bram[50633] = 219;
// bram[50634] = 234;
// bram[50635] = 245;
// bram[50636] = 252;
// bram[50637] = 253;
// bram[50638] = 251;
// bram[50639] = 243;
// bram[50640] = 232;
// bram[50641] = 216;
// bram[50642] = 197;
// bram[50643] = 175;
// bram[50644] = 152;
// bram[50645] = 127;
// bram[50646] = 103;
// bram[50647] = 79;
// bram[50648] = 57;
// bram[50649] = 38;
// bram[50650] = 22;
// bram[50651] = 10;
// bram[50652] = 3;
// bram[50653] = 0;
// bram[50654] = 1;
// bram[50655] = 8;
// bram[50656] = 18;
// bram[50657] = 33;
// bram[50658] = 52;
// bram[50659] = 73;
// bram[50660] = 96;
// bram[50661] = 120;
// bram[50662] = 145;
// bram[50663] = 169;
// bram[50664] = 191;
// bram[50665] = 211;
// bram[50666] = 227;
// bram[50667] = 240;
// bram[50668] = 249;
// bram[50669] = 253;
// bram[50670] = 253;
// bram[50671] = 247;
// bram[50672] = 237;
// bram[50673] = 223;
// bram[50674] = 206;
// bram[50675] = 185;
// bram[50676] = 163;
// bram[50677] = 138;
// bram[50678] = 114;
// bram[50679] = 90;
// bram[50680] = 67;
// bram[50681] = 47;
// bram[50682] = 29;
// bram[50683] = 15;
// bram[50684] = 6;
// bram[50685] = 0;
// bram[50686] = 0;
// bram[50687] = 4;
// bram[50688] = 13;
// bram[50689] = 26;
// bram[50690] = 43;
// bram[50691] = 63;
// bram[50692] = 85;
// bram[50693] = 109;
// bram[50694] = 134;
// bram[50695] = 158;
// bram[50696] = 181;
// bram[50697] = 202;
// bram[50698] = 220;
// bram[50699] = 235;
// bram[50700] = 246;
// bram[50701] = 252;
// bram[50702] = 253;
// bram[50703] = 250;
// bram[50704] = 242;
// bram[50705] = 230;
// bram[50706] = 214;
// bram[50707] = 195;
// bram[50708] = 173;
// bram[50709] = 149;
// bram[50710] = 125;
// bram[50711] = 101;
// bram[50712] = 77;
// bram[50713] = 56;
// bram[50714] = 37;
// bram[50715] = 21;
// bram[50716] = 9;
// bram[50717] = 2;
// bram[50718] = 0;
// bram[50719] = 2;
// bram[50720] = 8;
// bram[50721] = 20;
// bram[50722] = 35;
// bram[50723] = 53;
// bram[50724] = 75;
// bram[50725] = 98;
// bram[50726] = 122;
// bram[50727] = 147;
// bram[50728] = 171;
// bram[50729] = 193;
// bram[50730] = 212;
// bram[50731] = 229;
// bram[50732] = 241;
// bram[50733] = 250;
// bram[50734] = 253;
// bram[50735] = 252;
// bram[50736] = 247;
// bram[50737] = 236;
// bram[50738] = 222;
// bram[50739] = 204;
// bram[50740] = 183;
// bram[50741] = 160;
// bram[50742] = 136;
// bram[50743] = 112;
// bram[50744] = 88;
// bram[50745] = 65;
// bram[50746] = 45;
// bram[50747] = 28;
// bram[50748] = 14;
// bram[50749] = 5;
// bram[50750] = 0;
// bram[50751] = 0;
// bram[50752] = 5;
// bram[50753] = 14;
// bram[50754] = 27;
// bram[50755] = 45;
// bram[50756] = 65;
// bram[50757] = 87;
// bram[50758] = 111;
// bram[50759] = 136;
// bram[50760] = 160;
// bram[50761] = 183;
// bram[50762] = 204;
// bram[50763] = 222;
// bram[50764] = 236;
// bram[50765] = 246;
// bram[50766] = 252;
// bram[50767] = 253;
// bram[50768] = 250;
// bram[50769] = 241;
// bram[50770] = 229;
// bram[50771] = 213;
// bram[50772] = 193;
// bram[50773] = 171;
// bram[50774] = 147;
// bram[50775] = 123;
// bram[50776] = 98;
// bram[50777] = 75;
// bram[50778] = 54;
// bram[50779] = 35;
// bram[50780] = 20;
// bram[50781] = 9;
// bram[50782] = 2;
// bram[50783] = 0;
// bram[50784] = 2;
// bram[50785] = 9;
// bram[50786] = 21;
// bram[50787] = 36;
// bram[50788] = 55;
// bram[50789] = 77;
// bram[50790] = 100;
// bram[50791] = 125;
// bram[50792] = 149;
// bram[50793] = 173;
// bram[50794] = 195;
// bram[50795] = 214;
// bram[50796] = 230;
// bram[50797] = 242;
// bram[50798] = 250;
// bram[50799] = 253;
// bram[50800] = 252;
// bram[50801] = 246;
// bram[50802] = 235;
// bram[50803] = 220;
// bram[50804] = 202;
// bram[50805] = 181;
// bram[50806] = 158;
// bram[50807] = 134;
// bram[50808] = 109;
// bram[50809] = 86;
// bram[50810] = 63;
// bram[50811] = 43;
// bram[50812] = 26;
// bram[50813] = 13;
// bram[50814] = 4;
// bram[50815] = 0;
// bram[50816] = 0;
// bram[50817] = 5;
// bram[50818] = 15;
// bram[50819] = 29;
// bram[50820] = 46;
// bram[50821] = 67;
// bram[50822] = 89;
// bram[50823] = 114;
// bram[50824] = 138;
// bram[50825] = 162;
// bram[50826] = 185;
// bram[50827] = 206;
// bram[50828] = 223;
// bram[50829] = 237;
// bram[50830] = 247;
// bram[50831] = 253;
// bram[50832] = 253;
// bram[50833] = 249;
// bram[50834] = 241;
// bram[50835] = 228;
// bram[50836] = 211;
// bram[50837] = 191;
// bram[50838] = 169;
// bram[50839] = 145;
// bram[50840] = 121;
// bram[50841] = 96;
// bram[50842] = 73;
// bram[50843] = 52;
// bram[50844] = 34;
// bram[50845] = 19;
// bram[50846] = 8;
// bram[50847] = 1;
// bram[50848] = 0;
// bram[50849] = 3;
// bram[50850] = 10;
// bram[50851] = 22;
// bram[50852] = 38;
// bram[50853] = 57;
// bram[50854] = 79;
// bram[50855] = 102;
// bram[50856] = 127;
// bram[50857] = 151;
// bram[50858] = 175;
// bram[50859] = 197;
// bram[50860] = 216;
// bram[50861] = 231;
// bram[50862] = 243;
// bram[50863] = 251;
// bram[50864] = 253;
// bram[50865] = 252;
// bram[50866] = 245;
// bram[50867] = 234;
// bram[50868] = 219;
// bram[50869] = 200;
// bram[50870] = 179;
// bram[50871] = 156;
// bram[50872] = 132;
// bram[50873] = 107;
// bram[50874] = 83;
// bram[50875] = 61;
// bram[50876] = 41;
// bram[50877] = 25;
// bram[50878] = 12;
// bram[50879] = 4;
// bram[50880] = 0;
// bram[50881] = 1;
// bram[50882] = 6;
// bram[50883] = 16;
// bram[50884] = 30;
// bram[50885] = 48;
// bram[50886] = 69;
// bram[50887] = 92;
// bram[50888] = 116;
// bram[50889] = 140;
// bram[50890] = 164;
// bram[50891] = 187;
// bram[50892] = 207;
// bram[50893] = 225;
// bram[50894] = 238;
// bram[50895] = 248;
// bram[50896] = 253;
// bram[50897] = 253;
// bram[50898] = 249;
// bram[50899] = 239;
// bram[50900] = 226;
// bram[50901] = 209;
// bram[50902] = 189;
// bram[50903] = 167;
// bram[50904] = 143;
// bram[50905] = 118;
// bram[50906] = 94;
// bram[50907] = 71;
// bram[50908] = 50;
// bram[50909] = 32;
// bram[50910] = 17;
// bram[50911] = 7;
// bram[50912] = 1;
// bram[50913] = 0;
// bram[50914] = 3;
// bram[50915] = 11;
// bram[50916] = 23;
// bram[50917] = 40;
// bram[50918] = 59;
// bram[50919] = 81;
// bram[50920] = 105;
// bram[50921] = 129;
// bram[50922] = 154;
// bram[50923] = 177;
// bram[50924] = 198;
// bram[50925] = 217;
// bram[50926] = 233;
// bram[50927] = 244;
// bram[50928] = 251;
// bram[50929] = 253;
// bram[50930] = 251;
// bram[50931] = 244;
// bram[50932] = 233;
// bram[50933] = 217;
// bram[50934] = 199;
// bram[50935] = 177;
// bram[50936] = 154;
// bram[50937] = 129;
// bram[50938] = 105;
// bram[50939] = 81;
// bram[50940] = 59;
// bram[50941] = 40;
// bram[50942] = 24;
// bram[50943] = 11;
// bram[50944] = 3;
// bram[50945] = 0;
// bram[50946] = 1;
// bram[50947] = 7;
// bram[50948] = 17;
// bram[50949] = 32;
// bram[50950] = 50;
// bram[50951] = 71;
// bram[50952] = 94;
// bram[50953] = 118;
// bram[50954] = 143;
// bram[50955] = 166;
// bram[50956] = 189;
// bram[50957] = 209;
// bram[50958] = 226;
// bram[50959] = 239;
// bram[50960] = 248;
// bram[50961] = 253;
// bram[50962] = 253;
// bram[50963] = 248;
// bram[50964] = 238;
// bram[50965] = 225;
// bram[50966] = 208;
// bram[50967] = 187;
// bram[50968] = 165;
// bram[50969] = 141;
// bram[50970] = 116;
// bram[50971] = 92;
// bram[50972] = 69;
// bram[50973] = 48;
// bram[50974] = 31;
// bram[50975] = 16;
// bram[50976] = 6;
// bram[50977] = 1;
// bram[50978] = 0;
// bram[50979] = 4;
// bram[50980] = 12;
// bram[50981] = 25;
// bram[50982] = 41;
// bram[50983] = 61;
// bram[50984] = 83;
// bram[50985] = 107;
// bram[50986] = 131;
// bram[50987] = 156;
// bram[50988] = 179;
// bram[50989] = 200;
// bram[50990] = 219;
// bram[50991] = 234;
// bram[50992] = 245;
// bram[50993] = 252;
// bram[50994] = 253;
// bram[50995] = 251;
// bram[50996] = 243;
// bram[50997] = 232;
// bram[50998] = 216;
// bram[50999] = 197;
// bram[51000] = 175;
// bram[51001] = 152;
// bram[51002] = 127;
// bram[51003] = 103;
// bram[51004] = 79;
// bram[51005] = 57;
// bram[51006] = 38;
// bram[51007] = 22;
// bram[51008] = 10;
// bram[51009] = 3;
// bram[51010] = 0;
// bram[51011] = 1;
// bram[51012] = 8;
// bram[51013] = 18;
// bram[51014] = 33;
// bram[51015] = 52;
// bram[51016] = 73;
// bram[51017] = 96;
// bram[51018] = 120;
// bram[51019] = 145;
// bram[51020] = 169;
// bram[51021] = 191;
// bram[51022] = 211;
// bram[51023] = 227;
// bram[51024] = 240;
// bram[51025] = 249;
// bram[51026] = 253;
// bram[51027] = 253;
// bram[51028] = 247;
// bram[51029] = 237;
// bram[51030] = 223;
// bram[51031] = 206;
// bram[51032] = 185;
// bram[51033] = 162;
// bram[51034] = 138;
// bram[51035] = 114;
// bram[51036] = 90;
// bram[51037] = 67;
// bram[51038] = 47;
// bram[51039] = 29;
// bram[51040] = 15;
// bram[51041] = 6;
// bram[51042] = 0;
// bram[51043] = 0;
// bram[51044] = 4;
// bram[51045] = 13;
// bram[51046] = 26;
// bram[51047] = 43;
// bram[51048] = 63;
// bram[51049] = 85;
// bram[51050] = 109;
// bram[51051] = 134;
// bram[51052] = 158;
// bram[51053] = 181;
// bram[51054] = 202;
// bram[51055] = 220;
// bram[51056] = 235;
// bram[51057] = 246;
// bram[51058] = 252;
// bram[51059] = 253;
// bram[51060] = 250;
// bram[51061] = 242;
// bram[51062] = 230;
// bram[51063] = 214;
// bram[51064] = 195;
// bram[51065] = 173;
// bram[51066] = 149;
// bram[51067] = 125;
// bram[51068] = 101;
// bram[51069] = 77;
// bram[51070] = 56;
// bram[51071] = 37;
// bram[51072] = 21;
// bram[51073] = 9;
// bram[51074] = 2;
// bram[51075] = 0;
// bram[51076] = 2;
// bram[51077] = 8;
// bram[51078] = 20;
// bram[51079] = 35;
// bram[51080] = 53;
// bram[51081] = 75;
// bram[51082] = 98;
// bram[51083] = 122;
// bram[51084] = 147;
// bram[51085] = 171;
// bram[51086] = 193;
// bram[51087] = 212;
// bram[51088] = 229;
// bram[51089] = 241;
// bram[51090] = 250;
// bram[51091] = 253;
// bram[51092] = 252;
// bram[51093] = 247;
// bram[51094] = 236;
// bram[51095] = 222;
// bram[51096] = 204;
// bram[51097] = 183;
// bram[51098] = 160;
// bram[51099] = 136;
// bram[51100] = 112;
// bram[51101] = 88;
// bram[51102] = 65;
// bram[51103] = 45;
// bram[51104] = 28;
// bram[51105] = 14;
// bram[51106] = 5;
// bram[51107] = 0;
// bram[51108] = 0;
// bram[51109] = 5;
// bram[51110] = 14;
// bram[51111] = 27;
// bram[51112] = 45;
// bram[51113] = 65;
// bram[51114] = 87;
// bram[51115] = 111;
// bram[51116] = 136;
// bram[51117] = 160;
// bram[51118] = 183;
// bram[51119] = 204;
// bram[51120] = 222;
// bram[51121] = 236;
// bram[51122] = 246;
// bram[51123] = 252;
// bram[51124] = 253;
// bram[51125] = 250;
// bram[51126] = 241;
// bram[51127] = 229;
// bram[51128] = 213;
// bram[51129] = 193;
// bram[51130] = 171;
// bram[51131] = 147;
// bram[51132] = 123;
// bram[51133] = 98;
// bram[51134] = 75;
// bram[51135] = 54;
// bram[51136] = 35;
// bram[51137] = 20;
// bram[51138] = 9;
// bram[51139] = 2;
// bram[51140] = 0;
// bram[51141] = 2;
// bram[51142] = 9;
// bram[51143] = 21;
// bram[51144] = 36;
// bram[51145] = 55;
// bram[51146] = 77;
// bram[51147] = 100;
// bram[51148] = 125;
// bram[51149] = 149;
// bram[51150] = 173;
// bram[51151] = 195;
// bram[51152] = 214;
// bram[51153] = 230;
// bram[51154] = 242;
// bram[51155] = 250;
// bram[51156] = 253;
// bram[51157] = 252;
// bram[51158] = 246;
// bram[51159] = 235;
// bram[51160] = 220;
// bram[51161] = 202;
// bram[51162] = 181;
// bram[51163] = 158;
// bram[51164] = 134;
// bram[51165] = 109;
// bram[51166] = 85;
// bram[51167] = 63;
// bram[51168] = 43;
// bram[51169] = 26;
// bram[51170] = 13;
// bram[51171] = 4;
// bram[51172] = 0;
// bram[51173] = 0;
// bram[51174] = 5;
// bram[51175] = 15;
// bram[51176] = 29;
// bram[51177] = 46;
// bram[51178] = 67;
// bram[51179] = 89;
// bram[51180] = 114;
// bram[51181] = 138;
// bram[51182] = 162;
// bram[51183] = 185;
// bram[51184] = 206;
// bram[51185] = 223;
// bram[51186] = 237;
// bram[51187] = 247;
// bram[51188] = 253;
// bram[51189] = 253;
// bram[51190] = 249;
// bram[51191] = 240;
// bram[51192] = 228;
// bram[51193] = 211;
// bram[51194] = 191;
// bram[51195] = 169;
// bram[51196] = 145;
// bram[51197] = 120;
// bram[51198] = 96;
// bram[51199] = 73;
// bram[51200] = 52;
// bram[51201] = 33;
// bram[51202] = 19;
// bram[51203] = 8;
// bram[51204] = 1;
// bram[51205] = 0;
// bram[51206] = 3;
// bram[51207] = 10;
// bram[51208] = 22;
// bram[51209] = 38;
// bram[51210] = 57;
// bram[51211] = 79;
// bram[51212] = 103;
// bram[51213] = 127;
// bram[51214] = 151;
// bram[51215] = 175;
// bram[51216] = 197;
// bram[51217] = 216;
// bram[51218] = 231;
// bram[51219] = 243;
// bram[51220] = 251;
// bram[51221] = 253;
// bram[51222] = 252;
// bram[51223] = 245;
// bram[51224] = 234;
// bram[51225] = 219;
// bram[51226] = 200;
// bram[51227] = 179;
// bram[51228] = 156;
// bram[51229] = 132;
// bram[51230] = 107;
// bram[51231] = 83;
// bram[51232] = 61;
// bram[51233] = 41;
// bram[51234] = 25;
// bram[51235] = 12;
// bram[51236] = 4;
// bram[51237] = 0;
// bram[51238] = 1;
// bram[51239] = 6;
// bram[51240] = 16;
// bram[51241] = 30;
// bram[51242] = 48;
// bram[51243] = 69;
// bram[51244] = 92;
// bram[51245] = 116;
// bram[51246] = 140;
// bram[51247] = 164;
// bram[51248] = 187;
// bram[51249] = 207;
// bram[51250] = 225;
// bram[51251] = 238;
// bram[51252] = 248;
// bram[51253] = 253;
// bram[51254] = 253;
// bram[51255] = 249;
// bram[51256] = 239;
// bram[51257] = 226;
// bram[51258] = 209;
// bram[51259] = 189;
// bram[51260] = 167;
// bram[51261] = 143;
// bram[51262] = 118;
// bram[51263] = 94;
// bram[51264] = 71;
// bram[51265] = 50;
// bram[51266] = 32;
// bram[51267] = 17;
// bram[51268] = 7;
// bram[51269] = 1;
// bram[51270] = 0;
// bram[51271] = 3;
// bram[51272] = 11;
// bram[51273] = 23;
// bram[51274] = 40;
// bram[51275] = 59;
// bram[51276] = 81;
// bram[51277] = 105;
// bram[51278] = 129;
// bram[51279] = 154;
// bram[51280] = 177;
// bram[51281] = 198;
// bram[51282] = 217;
// bram[51283] = 233;
// bram[51284] = 244;
// bram[51285] = 251;
// bram[51286] = 253;
// bram[51287] = 251;
// bram[51288] = 244;
// bram[51289] = 233;
// bram[51290] = 217;
// bram[51291] = 199;
// bram[51292] = 177;
// bram[51293] = 154;
// bram[51294] = 129;
// bram[51295] = 105;
// bram[51296] = 81;
// bram[51297] = 59;
// bram[51298] = 40;
// bram[51299] = 24;
// bram[51300] = 11;
// bram[51301] = 3;
// bram[51302] = 0;
// bram[51303] = 1;
// bram[51304] = 7;
// bram[51305] = 17;
// bram[51306] = 32;
// bram[51307] = 50;
// bram[51308] = 71;
// bram[51309] = 94;
// bram[51310] = 118;
// bram[51311] = 143;
// bram[51312] = 167;
// bram[51313] = 189;
// bram[51314] = 209;
// bram[51315] = 226;
// bram[51316] = 239;
// bram[51317] = 248;
// bram[51318] = 253;
// bram[51319] = 253;
// bram[51320] = 248;
// bram[51321] = 238;
// bram[51322] = 225;
// bram[51323] = 207;
// bram[51324] = 187;
// bram[51325] = 165;
// bram[51326] = 141;
// bram[51327] = 116;
// bram[51328] = 92;
// bram[51329] = 69;
// bram[51330] = 48;
// bram[51331] = 30;
// bram[51332] = 16;
// bram[51333] = 6;
// bram[51334] = 1;
// bram[51335] = 0;
// bram[51336] = 4;
// bram[51337] = 12;
// bram[51338] = 25;
// bram[51339] = 41;
// bram[51340] = 61;
// bram[51341] = 83;
// bram[51342] = 107;
// bram[51343] = 131;
// bram[51344] = 156;
// bram[51345] = 179;
// bram[51346] = 200;
// bram[51347] = 219;
// bram[51348] = 234;
// bram[51349] = 245;
// bram[51350] = 252;
// bram[51351] = 253;
// bram[51352] = 251;
// bram[51353] = 243;
// bram[51354] = 231;
// bram[51355] = 216;
// bram[51356] = 197;
// bram[51357] = 175;
// bram[51358] = 152;
// bram[51359] = 127;
// bram[51360] = 103;
// bram[51361] = 79;
// bram[51362] = 57;
// bram[51363] = 38;
// bram[51364] = 22;
// bram[51365] = 10;
// bram[51366] = 3;
// bram[51367] = 0;
// bram[51368] = 1;
// bram[51369] = 8;
// bram[51370] = 18;
// bram[51371] = 33;
// bram[51372] = 52;
// bram[51373] = 73;
// bram[51374] = 96;
// bram[51375] = 120;
// bram[51376] = 145;
// bram[51377] = 169;
// bram[51378] = 191;
// bram[51379] = 211;
// bram[51380] = 227;
// bram[51381] = 240;
// bram[51382] = 249;
// bram[51383] = 253;
// bram[51384] = 253;
// bram[51385] = 247;
// bram[51386] = 237;
// bram[51387] = 223;
// bram[51388] = 206;
// bram[51389] = 185;
// bram[51390] = 162;
// bram[51391] = 138;
// bram[51392] = 114;
// bram[51393] = 90;
// bram[51394] = 67;
// bram[51395] = 47;
// bram[51396] = 29;
// bram[51397] = 15;
// bram[51398] = 6;
// bram[51399] = 0;
// bram[51400] = 0;
// bram[51401] = 4;
// bram[51402] = 13;
// bram[51403] = 26;
// bram[51404] = 43;
// bram[51405] = 63;
// bram[51406] = 85;
// bram[51407] = 109;
// bram[51408] = 134;
// bram[51409] = 158;
// bram[51410] = 181;
// bram[51411] = 202;
// bram[51412] = 220;
// bram[51413] = 235;
// bram[51414] = 246;
// bram[51415] = 252;
// bram[51416] = 253;
// bram[51417] = 250;
// bram[51418] = 242;
// bram[51419] = 230;
// bram[51420] = 214;
// bram[51421] = 195;
// bram[51422] = 173;
// bram[51423] = 149;
// bram[51424] = 125;
// bram[51425] = 101;
// bram[51426] = 77;
// bram[51427] = 55;
// bram[51428] = 37;
// bram[51429] = 21;
// bram[51430] = 9;
// bram[51431] = 2;
// bram[51432] = 0;
// bram[51433] = 2;
// bram[51434] = 8;
// bram[51435] = 20;
// bram[51436] = 35;
// bram[51437] = 54;
// bram[51438] = 75;
// bram[51439] = 98;
// bram[51440] = 123;
// bram[51441] = 147;
// bram[51442] = 171;
// bram[51443] = 193;
// bram[51444] = 212;
// bram[51445] = 229;
// bram[51446] = 241;
// bram[51447] = 250;
// bram[51448] = 253;
// bram[51449] = 252;
// bram[51450] = 246;
// bram[51451] = 236;
// bram[51452] = 222;
// bram[51453] = 204;
// bram[51454] = 183;
// bram[51455] = 160;
// bram[51456] = 136;
// bram[51457] = 112;
// bram[51458] = 88;
// bram[51459] = 65;
// bram[51460] = 45;
// bram[51461] = 28;
// bram[51462] = 14;
// bram[51463] = 5;
// bram[51464] = 0;
// bram[51465] = 0;
// bram[51466] = 5;
// bram[51467] = 14;
// bram[51468] = 28;
// bram[51469] = 45;
// bram[51470] = 65;
// bram[51471] = 87;
// bram[51472] = 111;
// bram[51473] = 136;
// bram[51474] = 160;
// bram[51475] = 183;
// bram[51476] = 204;
// bram[51477] = 222;
// bram[51478] = 236;
// bram[51479] = 246;
// bram[51480] = 252;
// bram[51481] = 253;
// bram[51482] = 250;
// bram[51483] = 241;
// bram[51484] = 229;
// bram[51485] = 213;
// bram[51486] = 193;
// bram[51487] = 171;
// bram[51488] = 147;
// bram[51489] = 123;
// bram[51490] = 98;
// bram[51491] = 75;
// bram[51492] = 54;
// bram[51493] = 35;
// bram[51494] = 20;
// bram[51495] = 9;
// bram[51496] = 2;
// bram[51497] = 0;
// bram[51498] = 2;
// bram[51499] = 9;
// bram[51500] = 21;
// bram[51501] = 36;
// bram[51502] = 55;
// bram[51503] = 77;
// bram[51504] = 100;
// bram[51505] = 125;
// bram[51506] = 149;
// bram[51507] = 173;
// bram[51508] = 195;
// bram[51509] = 214;
// bram[51510] = 230;
// bram[51511] = 242;
// bram[51512] = 250;
// bram[51513] = 253;
// bram[51514] = 252;
// bram[51515] = 246;
// bram[51516] = 235;
// bram[51517] = 220;
// bram[51518] = 202;
// bram[51519] = 181;
// bram[51520] = 158;
// bram[51521] = 134;
// bram[51522] = 109;
// bram[51523] = 85;
// bram[51524] = 63;
// bram[51525] = 43;
// bram[51526] = 26;
// bram[51527] = 13;
// bram[51528] = 4;
// bram[51529] = 0;
// bram[51530] = 0;
// bram[51531] = 5;
// bram[51532] = 15;
// bram[51533] = 29;
// bram[51534] = 46;
// bram[51535] = 67;
// bram[51536] = 90;
// bram[51537] = 114;
// bram[51538] = 138;
// bram[51539] = 162;
// bram[51540] = 185;
// bram[51541] = 206;
// bram[51542] = 223;
// bram[51543] = 237;
// bram[51544] = 247;
// bram[51545] = 253;
// bram[51546] = 253;
// bram[51547] = 249;
// bram[51548] = 240;
// bram[51549] = 228;
// bram[51550] = 211;
// bram[51551] = 191;
// bram[51552] = 169;
// bram[51553] = 145;
// bram[51554] = 120;
// bram[51555] = 96;
// bram[51556] = 73;
// bram[51557] = 52;
// bram[51558] = 33;
// bram[51559] = 19;
// bram[51560] = 8;
// bram[51561] = 1;
// bram[51562] = 0;
// bram[51563] = 3;
// bram[51564] = 10;
// bram[51565] = 22;
// bram[51566] = 38;
// bram[51567] = 57;
// bram[51568] = 79;
// bram[51569] = 103;
// bram[51570] = 127;
// bram[51571] = 151;
// bram[51572] = 175;
// bram[51573] = 197;
// bram[51574] = 216;
// bram[51575] = 231;
// bram[51576] = 243;
// bram[51577] = 251;
// bram[51578] = 253;
// bram[51579] = 252;
// bram[51580] = 245;
// bram[51581] = 234;
// bram[51582] = 219;
// bram[51583] = 200;
// bram[51584] = 179;
// bram[51585] = 156;
// bram[51586] = 132;
// bram[51587] = 107;
// bram[51588] = 83;
// bram[51589] = 61;
// bram[51590] = 41;
// bram[51591] = 25;
// bram[51592] = 12;
// bram[51593] = 4;
// bram[51594] = 0;
// bram[51595] = 1;
// bram[51596] = 6;
// bram[51597] = 16;
// bram[51598] = 30;
// bram[51599] = 48;
// bram[51600] = 69;
// bram[51601] = 92;
// bram[51602] = 116;
// bram[51603] = 140;
// bram[51604] = 164;
// bram[51605] = 187;
// bram[51606] = 207;
// bram[51607] = 225;
// bram[51608] = 238;
// bram[51609] = 248;
// bram[51610] = 253;
// bram[51611] = 253;
// bram[51612] = 249;
// bram[51613] = 239;
// bram[51614] = 226;
// bram[51615] = 209;
// bram[51616] = 189;
// bram[51617] = 167;
// bram[51618] = 143;
// bram[51619] = 118;
// bram[51620] = 94;
// bram[51621] = 71;
// bram[51622] = 50;
// bram[51623] = 32;
// bram[51624] = 17;
// bram[51625] = 7;
// bram[51626] = 1;
// bram[51627] = 0;
// bram[51628] = 3;
// bram[51629] = 11;
// bram[51630] = 23;
// bram[51631] = 40;
// bram[51632] = 59;
// bram[51633] = 81;
// bram[51634] = 105;
// bram[51635] = 129;
// bram[51636] = 154;
// bram[51637] = 177;
// bram[51638] = 198;
// bram[51639] = 217;
// bram[51640] = 233;
// bram[51641] = 244;
// bram[51642] = 251;
// bram[51643] = 253;
// bram[51644] = 251;
// bram[51645] = 244;
// bram[51646] = 233;
// bram[51647] = 217;
// bram[51648] = 199;
// bram[51649] = 177;
// bram[51650] = 154;
// bram[51651] = 129;
// bram[51652] = 105;
// bram[51653] = 81;
// bram[51654] = 59;
// bram[51655] = 40;
// bram[51656] = 24;
// bram[51657] = 11;
// bram[51658] = 3;
// bram[51659] = 0;
// bram[51660] = 1;
// bram[51661] = 7;
// bram[51662] = 17;
// bram[51663] = 32;
// bram[51664] = 50;
// bram[51665] = 71;
// bram[51666] = 94;
// bram[51667] = 118;
// bram[51668] = 143;
// bram[51669] = 167;
// bram[51670] = 189;
// bram[51671] = 209;
// bram[51672] = 226;
// bram[51673] = 239;
// bram[51674] = 248;
// bram[51675] = 253;
// bram[51676] = 253;
// bram[51677] = 248;
// bram[51678] = 238;
// bram[51679] = 225;
// bram[51680] = 207;
// bram[51681] = 187;
// bram[51682] = 165;
// bram[51683] = 140;
// bram[51684] = 116;
// bram[51685] = 92;
// bram[51686] = 69;
// bram[51687] = 48;
// bram[51688] = 30;
// bram[51689] = 16;
// bram[51690] = 6;
// bram[51691] = 1;
// bram[51692] = 0;
// bram[51693] = 4;
// bram[51694] = 12;
// bram[51695] = 25;
// bram[51696] = 41;
// bram[51697] = 61;
// bram[51698] = 83;
// bram[51699] = 107;
// bram[51700] = 131;
// bram[51701] = 156;
// bram[51702] = 179;
// bram[51703] = 200;
// bram[51704] = 219;
// bram[51705] = 234;
// bram[51706] = 245;
// bram[51707] = 252;
// bram[51708] = 253;
// bram[51709] = 251;
// bram[51710] = 243;
// bram[51711] = 231;
// bram[51712] = 216;
// bram[51713] = 197;
// bram[51714] = 175;
// bram[51715] = 152;
// bram[51716] = 127;
// bram[51717] = 103;
// bram[51718] = 79;
// bram[51719] = 57;
// bram[51720] = 38;
// bram[51721] = 22;
// bram[51722] = 10;
// bram[51723] = 3;
// bram[51724] = 0;
// bram[51725] = 1;
// bram[51726] = 8;
// bram[51727] = 19;
// bram[51728] = 33;
// bram[51729] = 52;
// bram[51730] = 73;
// bram[51731] = 96;
// bram[51732] = 120;
// bram[51733] = 145;
// bram[51734] = 169;
// bram[51735] = 191;
// bram[51736] = 211;
// bram[51737] = 227;
// bram[51738] = 240;
// bram[51739] = 249;
// bram[51740] = 253;
// bram[51741] = 253;
// bram[51742] = 247;
// bram[51743] = 237;
// bram[51744] = 223;
// bram[51745] = 206;
// bram[51746] = 185;
// bram[51747] = 162;
// bram[51748] = 138;
// bram[51749] = 114;
// bram[51750] = 90;
// bram[51751] = 67;
// bram[51752] = 46;
// bram[51753] = 29;
// bram[51754] = 15;
// bram[51755] = 5;
// bram[51756] = 0;
// bram[51757] = 0;
// bram[51758] = 4;
// bram[51759] = 13;
// bram[51760] = 26;
// bram[51761] = 43;
// bram[51762] = 63;
// bram[51763] = 85;
// bram[51764] = 109;
// bram[51765] = 134;
// bram[51766] = 158;
// bram[51767] = 181;
// bram[51768] = 202;
// bram[51769] = 220;
// bram[51770] = 235;
// bram[51771] = 246;
// bram[51772] = 252;
// bram[51773] = 253;
// bram[51774] = 250;
// bram[51775] = 242;
// bram[51776] = 230;
// bram[51777] = 214;
// bram[51778] = 195;
// bram[51779] = 173;
// bram[51780] = 149;
// bram[51781] = 125;
// bram[51782] = 100;
// bram[51783] = 77;
// bram[51784] = 55;
// bram[51785] = 37;
// bram[51786] = 21;
// bram[51787] = 9;
// bram[51788] = 2;
// bram[51789] = 0;
// bram[51790] = 2;
// bram[51791] = 8;
// bram[51792] = 20;
// bram[51793] = 35;
// bram[51794] = 54;
// bram[51795] = 75;
// bram[51796] = 98;
// bram[51797] = 123;
// bram[51798] = 147;
// bram[51799] = 171;
// bram[51800] = 193;
// bram[51801] = 212;
// bram[51802] = 229;
// bram[51803] = 241;
// bram[51804] = 250;
// bram[51805] = 253;
// bram[51806] = 252;
// bram[51807] = 246;
// bram[51808] = 236;
// bram[51809] = 222;
// bram[51810] = 204;
// bram[51811] = 183;
// bram[51812] = 160;
// bram[51813] = 136;
// bram[51814] = 111;
// bram[51815] = 87;
// bram[51816] = 65;
// bram[51817] = 45;
// bram[51818] = 28;
// bram[51819] = 14;
// bram[51820] = 5;
// bram[51821] = 0;
// bram[51822] = 0;
// bram[51823] = 5;
// bram[51824] = 14;
// bram[51825] = 28;
// bram[51826] = 45;
// bram[51827] = 65;
// bram[51828] = 87;
// bram[51829] = 111;
// bram[51830] = 136;
// bram[51831] = 160;
// bram[51832] = 183;
// bram[51833] = 204;
// bram[51834] = 222;
// bram[51835] = 236;
// bram[51836] = 246;
// bram[51837] = 252;
// bram[51838] = 253;
// bram[51839] = 250;
// bram[51840] = 241;
// bram[51841] = 229;
// bram[51842] = 212;
// bram[51843] = 193;
// bram[51844] = 171;
// bram[51845] = 147;
// bram[51846] = 123;
// bram[51847] = 98;
// bram[51848] = 75;
// bram[51849] = 54;
// bram[51850] = 35;
// bram[51851] = 20;
// bram[51852] = 8;
// bram[51853] = 2;
// bram[51854] = 0;
// bram[51855] = 2;
// bram[51856] = 9;
// bram[51857] = 21;
// bram[51858] = 36;
// bram[51859] = 55;
// bram[51860] = 77;
// bram[51861] = 100;
// bram[51862] = 125;
// bram[51863] = 149;
// bram[51864] = 173;
// bram[51865] = 195;
// bram[51866] = 214;
// bram[51867] = 230;
// bram[51868] = 242;
// bram[51869] = 250;
// bram[51870] = 253;
// bram[51871] = 252;
// bram[51872] = 246;
// bram[51873] = 235;
// bram[51874] = 220;
// bram[51875] = 202;
// bram[51876] = 181;
// bram[51877] = 158;
// bram[51878] = 134;
// bram[51879] = 109;
// bram[51880] = 85;
// bram[51881] = 63;
// bram[51882] = 43;
// bram[51883] = 26;
// bram[51884] = 13;
// bram[51885] = 4;
// bram[51886] = 0;
// bram[51887] = 0;
// bram[51888] = 5;
// bram[51889] = 15;
// bram[51890] = 29;
// bram[51891] = 46;
// bram[51892] = 67;
// bram[51893] = 90;
// bram[51894] = 114;
// bram[51895] = 138;
// bram[51896] = 162;
// bram[51897] = 185;
// bram[51898] = 206;
// bram[51899] = 223;
// bram[51900] = 237;
// bram[51901] = 247;
// bram[51902] = 253;
// bram[51903] = 253;
// bram[51904] = 249;
// bram[51905] = 240;
// bram[51906] = 228;
// bram[51907] = 211;
// bram[51908] = 191;
// bram[51909] = 169;
// bram[51910] = 145;
// bram[51911] = 120;
// bram[51912] = 96;
// bram[51913] = 73;
// bram[51914] = 52;
// bram[51915] = 33;
// bram[51916] = 19;
// bram[51917] = 8;
// bram[51918] = 1;
// bram[51919] = 0;
// bram[51920] = 3;
// bram[51921] = 10;
// bram[51922] = 22;
// bram[51923] = 38;
// bram[51924] = 57;
// bram[51925] = 79;
// bram[51926] = 103;
// bram[51927] = 127;
// bram[51928] = 151;
// bram[51929] = 175;
// bram[51930] = 197;
// bram[51931] = 216;
// bram[51932] = 231;
// bram[51933] = 243;
// bram[51934] = 251;
// bram[51935] = 253;
// bram[51936] = 252;
// bram[51937] = 245;
// bram[51938] = 234;
// bram[51939] = 219;
// bram[51940] = 200;
// bram[51941] = 179;
// bram[51942] = 156;
// bram[51943] = 132;
// bram[51944] = 107;
// bram[51945] = 83;
// bram[51946] = 61;
// bram[51947] = 41;
// bram[51948] = 25;
// bram[51949] = 12;
// bram[51950] = 4;
// bram[51951] = 0;
// bram[51952] = 1;
// bram[51953] = 6;
// bram[51954] = 16;
// bram[51955] = 30;
// bram[51956] = 48;
// bram[51957] = 69;
// bram[51958] = 92;
// bram[51959] = 116;
// bram[51960] = 140;
// bram[51961] = 164;
// bram[51962] = 187;
// bram[51963] = 207;
// bram[51964] = 225;
// bram[51965] = 238;
// bram[51966] = 248;
// bram[51967] = 253;
// bram[51968] = 253;
// bram[51969] = 248;
// bram[51970] = 239;
// bram[51971] = 226;
// bram[51972] = 209;
// bram[51973] = 189;
// bram[51974] = 167;
// bram[51975] = 143;
// bram[51976] = 118;
// bram[51977] = 94;
// bram[51978] = 71;
// bram[51979] = 50;
// bram[51980] = 32;
// bram[51981] = 17;
// bram[51982] = 7;
// bram[51983] = 1;
// bram[51984] = 0;
// bram[51985] = 3;
// bram[51986] = 11;
// bram[51987] = 23;
// bram[51988] = 40;
// bram[51989] = 59;
// bram[51990] = 81;
// bram[51991] = 105;
// bram[51992] = 129;
// bram[51993] = 154;
// bram[51994] = 177;
// bram[51995] = 199;
// bram[51996] = 217;
// bram[51997] = 233;
// bram[51998] = 244;
// bram[51999] = 251;
// bram[52000] = 254;
// bram[52001] = 251;
// bram[52002] = 244;
// bram[52003] = 233;
// bram[52004] = 217;
// bram[52005] = 199;
// bram[52006] = 177;
// bram[52007] = 154;
// bram[52008] = 129;
// bram[52009] = 105;
// bram[52010] = 81;
// bram[52011] = 59;
// bram[52012] = 40;
// bram[52013] = 23;
// bram[52014] = 11;
// bram[52015] = 3;
// bram[52016] = 0;
// bram[52017] = 1;
// bram[52018] = 7;
// bram[52019] = 17;
// bram[52020] = 32;
// bram[52021] = 50;
// bram[52022] = 71;
// bram[52023] = 94;
// bram[52024] = 118;
// bram[52025] = 143;
// bram[52026] = 167;
// bram[52027] = 189;
// bram[52028] = 209;
// bram[52029] = 226;
// bram[52030] = 239;
// bram[52031] = 248;
// bram[52032] = 253;
// bram[52033] = 253;
// bram[52034] = 248;
// bram[52035] = 238;
// bram[52036] = 225;
// bram[52037] = 207;
// bram[52038] = 187;
// bram[52039] = 164;
// bram[52040] = 140;
// bram[52041] = 116;
// bram[52042] = 92;
// bram[52043] = 69;
// bram[52044] = 48;
// bram[52045] = 30;
// bram[52046] = 16;
// bram[52047] = 6;
// bram[52048] = 1;
// bram[52049] = 0;
// bram[52050] = 4;
// bram[52051] = 12;
// bram[52052] = 25;
// bram[52053] = 41;
// bram[52054] = 61;
// bram[52055] = 83;
// bram[52056] = 107;
// bram[52057] = 132;
// bram[52058] = 156;
// bram[52059] = 179;
// bram[52060] = 200;
// bram[52061] = 219;
// bram[52062] = 234;
// bram[52063] = 245;
// bram[52064] = 252;
// bram[52065] = 253;
// bram[52066] = 251;
// bram[52067] = 243;
// bram[52068] = 231;
// bram[52069] = 216;
// bram[52070] = 197;
// bram[52071] = 175;
// bram[52072] = 151;
// bram[52073] = 127;
// bram[52074] = 103;
// bram[52075] = 79;
// bram[52076] = 57;
// bram[52077] = 38;
// bram[52078] = 22;
// bram[52079] = 10;
// bram[52080] = 3;
// bram[52081] = 0;
// bram[52082] = 1;
// bram[52083] = 8;
// bram[52084] = 19;
// bram[52085] = 33;
// bram[52086] = 52;
// bram[52087] = 73;
// bram[52088] = 96;
// bram[52089] = 120;
// bram[52090] = 145;
// bram[52091] = 169;
// bram[52092] = 191;
// bram[52093] = 211;
// bram[52094] = 228;
// bram[52095] = 240;
// bram[52096] = 249;
// bram[52097] = 253;
// bram[52098] = 253;
// bram[52099] = 247;
// bram[52100] = 237;
// bram[52101] = 223;
// bram[52102] = 206;
// bram[52103] = 185;
// bram[52104] = 162;
// bram[52105] = 138;
// bram[52106] = 114;
// bram[52107] = 90;
// bram[52108] = 67;
// bram[52109] = 46;
// bram[52110] = 29;
// bram[52111] = 15;
// bram[52112] = 5;
// bram[52113] = 0;
// bram[52114] = 0;
// bram[52115] = 4;
// bram[52116] = 13;
// bram[52117] = 26;
// bram[52118] = 43;
// bram[52119] = 63;
// bram[52120] = 85;
// bram[52121] = 109;
// bram[52122] = 134;
// bram[52123] = 158;
// bram[52124] = 181;
// bram[52125] = 202;
// bram[52126] = 220;
// bram[52127] = 235;
// bram[52128] = 246;
// bram[52129] = 252;
// bram[52130] = 253;
// bram[52131] = 250;
// bram[52132] = 242;
// bram[52133] = 230;
// bram[52134] = 214;
// bram[52135] = 195;
// bram[52136] = 173;
// bram[52137] = 149;
// bram[52138] = 125;
// bram[52139] = 100;
// bram[52140] = 77;
// bram[52141] = 55;
// bram[52142] = 36;
// bram[52143] = 21;
// bram[52144] = 9;
// bram[52145] = 2;
// bram[52146] = 0;
// bram[52147] = 2;
// bram[52148] = 8;
// bram[52149] = 20;
// bram[52150] = 35;
// bram[52151] = 54;
// bram[52152] = 75;
// bram[52153] = 98;
// bram[52154] = 123;
// bram[52155] = 147;
// bram[52156] = 171;
// bram[52157] = 193;
// bram[52158] = 212;
// bram[52159] = 229;
// bram[52160] = 241;
// bram[52161] = 250;
// bram[52162] = 253;
// bram[52163] = 252;
// bram[52164] = 246;
// bram[52165] = 236;
// bram[52166] = 222;
// bram[52167] = 204;
// bram[52168] = 183;
// bram[52169] = 160;
// bram[52170] = 136;
// bram[52171] = 111;
// bram[52172] = 87;
// bram[52173] = 65;
// bram[52174] = 45;
// bram[52175] = 28;
// bram[52176] = 14;
// bram[52177] = 5;
// bram[52178] = 0;
// bram[52179] = 0;
// bram[52180] = 5;
// bram[52181] = 14;
// bram[52182] = 28;
// bram[52183] = 45;
// bram[52184] = 65;
// bram[52185] = 87;
// bram[52186] = 111;
// bram[52187] = 136;
// bram[52188] = 160;
// bram[52189] = 183;
// bram[52190] = 204;
// bram[52191] = 222;
// bram[52192] = 236;
// bram[52193] = 246;
// bram[52194] = 252;
// bram[52195] = 253;
// bram[52196] = 250;
// bram[52197] = 241;
// bram[52198] = 229;
// bram[52199] = 212;
// bram[52200] = 193;
// bram[52201] = 171;
// bram[52202] = 147;
// bram[52203] = 123;
// bram[52204] = 98;
// bram[52205] = 75;
// bram[52206] = 54;
// bram[52207] = 35;
// bram[52208] = 20;
// bram[52209] = 8;
// bram[52210] = 2;
// bram[52211] = 0;
// bram[52212] = 2;
// bram[52213] = 9;
// bram[52214] = 21;
// bram[52215] = 37;
// bram[52216] = 55;
// bram[52217] = 77;
// bram[52218] = 100;
// bram[52219] = 125;
// bram[52220] = 149;
// bram[52221] = 173;
// bram[52222] = 195;
// bram[52223] = 214;
// bram[52224] = 230;
// bram[52225] = 242;
// bram[52226] = 250;
// bram[52227] = 253;
// bram[52228] = 252;
// bram[52229] = 246;
// bram[52230] = 235;
// bram[52231] = 220;
// bram[52232] = 202;
// bram[52233] = 181;
// bram[52234] = 158;
// bram[52235] = 134;
// bram[52236] = 109;
// bram[52237] = 85;
// bram[52238] = 63;
// bram[52239] = 43;
// bram[52240] = 26;
// bram[52241] = 13;
// bram[52242] = 4;
// bram[52243] = 0;
// bram[52244] = 0;
// bram[52245] = 5;
// bram[52246] = 15;
// bram[52247] = 29;
// bram[52248] = 46;
// bram[52249] = 67;
// bram[52250] = 90;
// bram[52251] = 114;
// bram[52252] = 138;
// bram[52253] = 162;
// bram[52254] = 185;
// bram[52255] = 206;
// bram[52256] = 223;
// bram[52257] = 237;
// bram[52258] = 247;
// bram[52259] = 253;
// bram[52260] = 253;
// bram[52261] = 249;
// bram[52262] = 240;
// bram[52263] = 227;
// bram[52264] = 211;
// bram[52265] = 191;
// bram[52266] = 169;
// bram[52267] = 145;
// bram[52268] = 120;
// bram[52269] = 96;
// bram[52270] = 73;
// bram[52271] = 52;
// bram[52272] = 33;
// bram[52273] = 19;
// bram[52274] = 8;
// bram[52275] = 1;
// bram[52276] = 0;
// bram[52277] = 3;
// bram[52278] = 10;
// bram[52279] = 22;
// bram[52280] = 38;
// bram[52281] = 57;
// bram[52282] = 79;
// bram[52283] = 103;
// bram[52284] = 127;
// bram[52285] = 152;
// bram[52286] = 175;
// bram[52287] = 197;
// bram[52288] = 216;
// bram[52289] = 231;
// bram[52290] = 243;
// bram[52291] = 251;
// bram[52292] = 253;
// bram[52293] = 252;
// bram[52294] = 245;
// bram[52295] = 234;
// bram[52296] = 219;
// bram[52297] = 200;
// bram[52298] = 179;
// bram[52299] = 156;
// bram[52300] = 131;
// bram[52301] = 107;
// bram[52302] = 83;
// bram[52303] = 61;
// bram[52304] = 41;
// bram[52305] = 25;
// bram[52306] = 12;
// bram[52307] = 4;
// bram[52308] = 0;
// bram[52309] = 1;
// bram[52310] = 6;
// bram[52311] = 16;
// bram[52312] = 30;
// bram[52313] = 48;
// bram[52314] = 69;
// bram[52315] = 92;
// bram[52316] = 116;
// bram[52317] = 140;
// bram[52318] = 165;
// bram[52319] = 187;
// bram[52320] = 207;
// bram[52321] = 225;
// bram[52322] = 238;
// bram[52323] = 248;
// bram[52324] = 253;
// bram[52325] = 253;
// bram[52326] = 248;
// bram[52327] = 239;
// bram[52328] = 226;
// bram[52329] = 209;
// bram[52330] = 189;
// bram[52331] = 167;
// bram[52332] = 143;
// bram[52333] = 118;
// bram[52334] = 94;
// bram[52335] = 71;
// bram[52336] = 50;
// bram[52337] = 32;
// bram[52338] = 17;
// bram[52339] = 7;
// bram[52340] = 1;
// bram[52341] = 0;
// bram[52342] = 3;
// bram[52343] = 11;
// bram[52344] = 24;
// bram[52345] = 40;
// bram[52346] = 59;
// bram[52347] = 81;
// bram[52348] = 105;
// bram[52349] = 129;
// bram[52350] = 154;
// bram[52351] = 177;
// bram[52352] = 199;
// bram[52353] = 217;
// bram[52354] = 233;
// bram[52355] = 244;
// bram[52356] = 251;
// bram[52357] = 253;
// bram[52358] = 251;
// bram[52359] = 244;
// bram[52360] = 233;
// bram[52361] = 217;
// bram[52362] = 198;
// bram[52363] = 177;
// bram[52364] = 154;
// bram[52365] = 129;
// bram[52366] = 105;
// bram[52367] = 81;
// bram[52368] = 59;
// bram[52369] = 40;
// bram[52370] = 23;
// bram[52371] = 11;
// bram[52372] = 3;
// bram[52373] = 0;
// bram[52374] = 1;
// bram[52375] = 7;
// bram[52376] = 17;
// bram[52377] = 32;
// bram[52378] = 50;
// bram[52379] = 71;
// bram[52380] = 94;
// bram[52381] = 118;
// bram[52382] = 143;
// bram[52383] = 167;
// bram[52384] = 189;
// bram[52385] = 209;
// bram[52386] = 226;
// bram[52387] = 239;
// bram[52388] = 249;
// bram[52389] = 253;
// bram[52390] = 253;
// bram[52391] = 248;
// bram[52392] = 238;
// bram[52393] = 225;
// bram[52394] = 207;
// bram[52395] = 187;
// bram[52396] = 164;
// bram[52397] = 140;
// bram[52398] = 116;
// bram[52399] = 92;
// bram[52400] = 69;
// bram[52401] = 48;
// bram[52402] = 30;
// bram[52403] = 16;
// bram[52404] = 6;
// bram[52405] = 1;
// bram[52406] = 0;
// bram[52407] = 4;
// bram[52408] = 12;
// bram[52409] = 25;
// bram[52410] = 41;
// bram[52411] = 61;
// bram[52412] = 83;
// bram[52413] = 107;
// bram[52414] = 132;
// bram[52415] = 156;
// bram[52416] = 179;
// bram[52417] = 200;
// bram[52418] = 219;
// bram[52419] = 234;
// bram[52420] = 245;
// bram[52421] = 252;
// bram[52422] = 253;
// bram[52423] = 251;
// bram[52424] = 243;
// bram[52425] = 231;
// bram[52426] = 216;
// bram[52427] = 197;
// bram[52428] = 175;
// bram[52429] = 151;
// bram[52430] = 127;
// bram[52431] = 103;
// bram[52432] = 79;
// bram[52433] = 57;
// bram[52434] = 38;
// bram[52435] = 22;
// bram[52436] = 10;
// bram[52437] = 3;
// bram[52438] = 0;
// bram[52439] = 1;
// bram[52440] = 8;
// bram[52441] = 19;
// bram[52442] = 33;
// bram[52443] = 52;
// bram[52444] = 73;
// bram[52445] = 96;
// bram[52446] = 120;
// bram[52447] = 145;
// bram[52448] = 169;
// bram[52449] = 191;
// bram[52450] = 211;
// bram[52451] = 228;
// bram[52452] = 240;
// bram[52453] = 249;
// bram[52454] = 253;
// bram[52455] = 253;
// bram[52456] = 247;
// bram[52457] = 237;
// bram[52458] = 223;
// bram[52459] = 206;
// bram[52460] = 185;
// bram[52461] = 162;
// bram[52462] = 138;
// bram[52463] = 114;
// bram[52464] = 90;
// bram[52465] = 67;
// bram[52466] = 46;
// bram[52467] = 29;
// bram[52468] = 15;
// bram[52469] = 5;
// bram[52470] = 0;
// bram[52471] = 0;
// bram[52472] = 4;
// bram[52473] = 13;
// bram[52474] = 26;
// bram[52475] = 43;
// bram[52476] = 63;
// bram[52477] = 85;
// bram[52478] = 109;
// bram[52479] = 134;
// bram[52480] = 158;
// bram[52481] = 181;
// bram[52482] = 202;
// bram[52483] = 220;
// bram[52484] = 235;
// bram[52485] = 246;
// bram[52486] = 252;
// bram[52487] = 253;
// bram[52488] = 250;
// bram[52489] = 242;
// bram[52490] = 230;
// bram[52491] = 214;
// bram[52492] = 195;
// bram[52493] = 173;
// bram[52494] = 149;
// bram[52495] = 125;
// bram[52496] = 100;
// bram[52497] = 77;
// bram[52498] = 55;
// bram[52499] = 36;
// bram[52500] = 21;
// bram[52501] = 9;
// bram[52502] = 2;
// bram[52503] = 0;
// bram[52504] = 2;
// bram[52505] = 9;
// bram[52506] = 20;
// bram[52507] = 35;
// bram[52508] = 54;
// bram[52509] = 75;
// bram[52510] = 98;
// bram[52511] = 123;
// bram[52512] = 147;
// bram[52513] = 171;
// bram[52514] = 193;
// bram[52515] = 213;
// bram[52516] = 229;
// bram[52517] = 241;
// bram[52518] = 250;
// bram[52519] = 253;
// bram[52520] = 252;
// bram[52521] = 246;
// bram[52522] = 236;
// bram[52523] = 222;
// bram[52524] = 204;
// bram[52525] = 183;
// bram[52526] = 160;
// bram[52527] = 136;
// bram[52528] = 111;
// bram[52529] = 87;
// bram[52530] = 65;
// bram[52531] = 45;
// bram[52532] = 28;
// bram[52533] = 14;
// bram[52534] = 5;
// bram[52535] = 0;
// bram[52536] = 0;
// bram[52537] = 5;
// bram[52538] = 14;
// bram[52539] = 28;
// bram[52540] = 45;
// bram[52541] = 65;
// bram[52542] = 88;
// bram[52543] = 112;
// bram[52544] = 136;
// bram[52545] = 160;
// bram[52546] = 183;
// bram[52547] = 204;
// bram[52548] = 222;
// bram[52549] = 236;
// bram[52550] = 246;
// bram[52551] = 252;
// bram[52552] = 253;
// bram[52553] = 250;
// bram[52554] = 241;
// bram[52555] = 229;
// bram[52556] = 212;
// bram[52557] = 193;
// bram[52558] = 171;
// bram[52559] = 147;
// bram[52560] = 123;
// bram[52561] = 98;
// bram[52562] = 75;
// bram[52563] = 54;
// bram[52564] = 35;
// bram[52565] = 20;
// bram[52566] = 8;
// bram[52567] = 2;
// bram[52568] = 0;
// bram[52569] = 2;
// bram[52570] = 9;
// bram[52571] = 21;
// bram[52572] = 37;
// bram[52573] = 55;
// bram[52574] = 77;
// bram[52575] = 101;
// bram[52576] = 125;
// bram[52577] = 149;
// bram[52578] = 173;
// bram[52579] = 195;
// bram[52580] = 214;
// bram[52581] = 230;
// bram[52582] = 242;
// bram[52583] = 250;
// bram[52584] = 253;
// bram[52585] = 252;
// bram[52586] = 246;
// bram[52587] = 235;
// bram[52588] = 220;
// bram[52589] = 202;
// bram[52590] = 181;
// bram[52591] = 158;
// bram[52592] = 134;
// bram[52593] = 109;
// bram[52594] = 85;
// bram[52595] = 63;
// bram[52596] = 43;
// bram[52597] = 26;
// bram[52598] = 13;
// bram[52599] = 4;
// bram[52600] = 0;
// bram[52601] = 0;
// bram[52602] = 6;
// bram[52603] = 15;
// bram[52604] = 29;
// bram[52605] = 47;
// bram[52606] = 67;
// bram[52607] = 90;
// bram[52608] = 114;
// bram[52609] = 138;
// bram[52610] = 162;
// bram[52611] = 185;
// bram[52612] = 206;
// bram[52613] = 223;
// bram[52614] = 237;
// bram[52615] = 247;
// bram[52616] = 253;
// bram[52617] = 253;
// bram[52618] = 249;
// bram[52619] = 240;
// bram[52620] = 227;
// bram[52621] = 211;
// bram[52622] = 191;
// bram[52623] = 169;
// bram[52624] = 145;
// bram[52625] = 120;
// bram[52626] = 96;
// bram[52627] = 73;
// bram[52628] = 52;
// bram[52629] = 33;
// bram[52630] = 18;
// bram[52631] = 8;
// bram[52632] = 1;
// bram[52633] = 0;
// bram[52634] = 3;
// bram[52635] = 10;
// bram[52636] = 22;
// bram[52637] = 38;
// bram[52638] = 57;
// bram[52639] = 79;
// bram[52640] = 103;
// bram[52641] = 127;
// bram[52642] = 152;
// bram[52643] = 175;
// bram[52644] = 197;
// bram[52645] = 216;
// bram[52646] = 231;
// bram[52647] = 243;
// bram[52648] = 251;
// bram[52649] = 253;
// bram[52650] = 252;
// bram[52651] = 245;
// bram[52652] = 234;
// bram[52653] = 219;
// bram[52654] = 200;
// bram[52655] = 179;
// bram[52656] = 156;
// bram[52657] = 131;
// bram[52658] = 107;
// bram[52659] = 83;
// bram[52660] = 61;
// bram[52661] = 41;
// bram[52662] = 25;
// bram[52663] = 12;
// bram[52664] = 4;
// bram[52665] = 0;
// bram[52666] = 1;
// bram[52667] = 6;
// bram[52668] = 16;
// bram[52669] = 30;
// bram[52670] = 48;
// bram[52671] = 69;
// bram[52672] = 92;
// bram[52673] = 116;
// bram[52674] = 141;
// bram[52675] = 165;
// bram[52676] = 187;
// bram[52677] = 207;
// bram[52678] = 225;
// bram[52679] = 238;
// bram[52680] = 248;
// bram[52681] = 253;
// bram[52682] = 253;
// bram[52683] = 248;
// bram[52684] = 239;
// bram[52685] = 226;
// bram[52686] = 209;
// bram[52687] = 189;
// bram[52688] = 167;
// bram[52689] = 143;
// bram[52690] = 118;
// bram[52691] = 94;
// bram[52692] = 71;
// bram[52693] = 50;
// bram[52694] = 32;
// bram[52695] = 17;
// bram[52696] = 7;
// bram[52697] = 1;
// bram[52698] = 0;
// bram[52699] = 3;
// bram[52700] = 11;
// bram[52701] = 24;
// bram[52702] = 40;
// bram[52703] = 59;
// bram[52704] = 81;
// bram[52705] = 105;
// bram[52706] = 129;
// bram[52707] = 154;
// bram[52708] = 177;
// bram[52709] = 199;
// bram[52710] = 217;
// bram[52711] = 233;
// bram[52712] = 244;
// bram[52713] = 251;
// bram[52714] = 253;
// bram[52715] = 251;
// bram[52716] = 244;
// bram[52717] = 233;
// bram[52718] = 217;
// bram[52719] = 198;
// bram[52720] = 177;
// bram[52721] = 154;
// bram[52722] = 129;
// bram[52723] = 105;
// bram[52724] = 81;
// bram[52725] = 59;
// bram[52726] = 40;
// bram[52727] = 23;
// bram[52728] = 11;
// bram[52729] = 3;
// bram[52730] = 0;
// bram[52731] = 1;
// bram[52732] = 7;
// bram[52733] = 17;
// bram[52734] = 32;
// bram[52735] = 50;
// bram[52736] = 71;
// bram[52737] = 94;
// bram[52738] = 118;
// bram[52739] = 143;
// bram[52740] = 167;
// bram[52741] = 189;
// bram[52742] = 209;
// bram[52743] = 226;
// bram[52744] = 239;
// bram[52745] = 249;
// bram[52746] = 253;
// bram[52747] = 253;
// bram[52748] = 248;
// bram[52749] = 238;
// bram[52750] = 225;
// bram[52751] = 207;
// bram[52752] = 187;
// bram[52753] = 164;
// bram[52754] = 140;
// bram[52755] = 116;
// bram[52756] = 92;
// bram[52757] = 69;
// bram[52758] = 48;
// bram[52759] = 30;
// bram[52760] = 16;
// bram[52761] = 6;
// bram[52762] = 1;
// bram[52763] = 0;
// bram[52764] = 4;
// bram[52765] = 12;
// bram[52766] = 25;
// bram[52767] = 41;
// bram[52768] = 61;
// bram[52769] = 83;
// bram[52770] = 107;
// bram[52771] = 132;
// bram[52772] = 156;
// bram[52773] = 179;
// bram[52774] = 200;
// bram[52775] = 219;
// bram[52776] = 234;
// bram[52777] = 245;
// bram[52778] = 252;
// bram[52779] = 253;
// bram[52780] = 251;
// bram[52781] = 243;
// bram[52782] = 231;
// bram[52783] = 216;
// bram[52784] = 197;
// bram[52785] = 175;
// bram[52786] = 151;
// bram[52787] = 127;
// bram[52788] = 103;
// bram[52789] = 79;
// bram[52790] = 57;
// bram[52791] = 38;
// bram[52792] = 22;
// bram[52793] = 10;
// bram[52794] = 3;
// bram[52795] = 0;
// bram[52796] = 1;
// bram[52797] = 8;
// bram[52798] = 19;
// bram[52799] = 33;
// bram[52800] = 52;
// bram[52801] = 73;
// bram[52802] = 96;
// bram[52803] = 120;
// bram[52804] = 145;
// bram[52805] = 169;
// bram[52806] = 191;
// bram[52807] = 211;
// bram[52808] = 228;
// bram[52809] = 240;
// bram[52810] = 249;
// bram[52811] = 253;
// bram[52812] = 253;
// bram[52813] = 247;
// bram[52814] = 237;
// bram[52815] = 223;
// bram[52816] = 206;
// bram[52817] = 185;
// bram[52818] = 162;
// bram[52819] = 138;
// bram[52820] = 114;
// bram[52821] = 89;
// bram[52822] = 67;
// bram[52823] = 46;
// bram[52824] = 29;
// bram[52825] = 15;
// bram[52826] = 5;
// bram[52827] = 0;
// bram[52828] = 0;
// bram[52829] = 4;
// bram[52830] = 13;
// bram[52831] = 26;
// bram[52832] = 43;
// bram[52833] = 63;
// bram[52834] = 85;
// bram[52835] = 109;
// bram[52836] = 134;
// bram[52837] = 158;
// bram[52838] = 181;
// bram[52839] = 202;
// bram[52840] = 220;
// bram[52841] = 235;
// bram[52842] = 246;
// bram[52843] = 252;
// bram[52844] = 253;
// bram[52845] = 250;
// bram[52846] = 242;
// bram[52847] = 230;
// bram[52848] = 214;
// bram[52849] = 195;
// bram[52850] = 173;
// bram[52851] = 149;
// bram[52852] = 125;
// bram[52853] = 100;
// bram[52854] = 77;
// bram[52855] = 55;
// bram[52856] = 36;
// bram[52857] = 21;
// bram[52858] = 9;
// bram[52859] = 2;
// bram[52860] = 0;
// bram[52861] = 2;
// bram[52862] = 9;
// bram[52863] = 20;
// bram[52864] = 35;
// bram[52865] = 54;
// bram[52866] = 75;
// bram[52867] = 98;
// bram[52868] = 123;
// bram[52869] = 147;
// bram[52870] = 171;
// bram[52871] = 193;
// bram[52872] = 213;
// bram[52873] = 229;
// bram[52874] = 241;
// bram[52875] = 250;
// bram[52876] = 253;
// bram[52877] = 252;
// bram[52878] = 246;
// bram[52879] = 236;
// bram[52880] = 222;
// bram[52881] = 204;
// bram[52882] = 183;
// bram[52883] = 160;
// bram[52884] = 136;
// bram[52885] = 111;
// bram[52886] = 87;
// bram[52887] = 65;
// bram[52888] = 45;
// bram[52889] = 27;
// bram[52890] = 14;
// bram[52891] = 5;
// bram[52892] = 0;
// bram[52893] = 0;
// bram[52894] = 5;
// bram[52895] = 14;
// bram[52896] = 28;
// bram[52897] = 45;
// bram[52898] = 65;
// bram[52899] = 88;
// bram[52900] = 112;
// bram[52901] = 136;
// bram[52902] = 160;
// bram[52903] = 183;
// bram[52904] = 204;
// bram[52905] = 222;
// bram[52906] = 236;
// bram[52907] = 247;
// bram[52908] = 252;
// bram[52909] = 253;
// bram[52910] = 250;
// bram[52911] = 241;
// bram[52912] = 229;
// bram[52913] = 212;
// bram[52914] = 193;
// bram[52915] = 171;
// bram[52916] = 147;
// bram[52917] = 122;
// bram[52918] = 98;
// bram[52919] = 75;
// bram[52920] = 53;
// bram[52921] = 35;
// bram[52922] = 20;
// bram[52923] = 8;
// bram[52924] = 2;
// bram[52925] = 0;
// bram[52926] = 2;
// bram[52927] = 9;
// bram[52928] = 21;
// bram[52929] = 37;
// bram[52930] = 56;
// bram[52931] = 77;
// bram[52932] = 101;
// bram[52933] = 125;
// bram[52934] = 149;
// bram[52935] = 173;
// bram[52936] = 195;
// bram[52937] = 214;
// bram[52938] = 230;
// bram[52939] = 242;
// bram[52940] = 250;
// bram[52941] = 253;
// bram[52942] = 252;
// bram[52943] = 246;
// bram[52944] = 235;
// bram[52945] = 220;
// bram[52946] = 202;
// bram[52947] = 181;
// bram[52948] = 158;
// bram[52949] = 134;
// bram[52950] = 109;
// bram[52951] = 85;
// bram[52952] = 63;
// bram[52953] = 43;
// bram[52954] = 26;
// bram[52955] = 13;
// bram[52956] = 4;
// bram[52957] = 0;
// bram[52958] = 0;
// bram[52959] = 6;
// bram[52960] = 15;
// bram[52961] = 29;
// bram[52962] = 47;
// bram[52963] = 67;
// bram[52964] = 90;
// bram[52965] = 114;
// bram[52966] = 138;
// bram[52967] = 162;
// bram[52968] = 185;
// bram[52969] = 206;
// bram[52970] = 223;
// bram[52971] = 237;
// bram[52972] = 247;
// bram[52973] = 253;
// bram[52974] = 253;
// bram[52975] = 249;
// bram[52976] = 240;
// bram[52977] = 227;
// bram[52978] = 211;
// bram[52979] = 191;
// bram[52980] = 169;
// bram[52981] = 145;
// bram[52982] = 120;
// bram[52983] = 96;
// bram[52984] = 73;
// bram[52985] = 52;
// bram[52986] = 33;
// bram[52987] = 18;
// bram[52988] = 8;
// bram[52989] = 1;
// bram[52990] = 0;
// bram[52991] = 3;
// bram[52992] = 10;
// bram[52993] = 22;
// bram[52994] = 38;
// bram[52995] = 57;
// bram[52996] = 79;
// bram[52997] = 103;
// bram[52998] = 127;
// bram[52999] = 152;
// bram[53000] = 175;
// bram[53001] = 197;
// bram[53002] = 216;
// bram[53003] = 232;
// bram[53004] = 243;
// bram[53005] = 251;
// bram[53006] = 253;
// bram[53007] = 252;
// bram[53008] = 245;
// bram[53009] = 234;
// bram[53010] = 219;
// bram[53011] = 200;
// bram[53012] = 179;
// bram[53013] = 156;
// bram[53014] = 131;
// bram[53015] = 107;
// bram[53016] = 83;
// bram[53017] = 61;
// bram[53018] = 41;
// bram[53019] = 25;
// bram[53020] = 12;
// bram[53021] = 4;
// bram[53022] = 0;
// bram[53023] = 1;
// bram[53024] = 6;
// bram[53025] = 16;
// bram[53026] = 31;
// bram[53027] = 48;
// bram[53028] = 69;
// bram[53029] = 92;
// bram[53030] = 116;
// bram[53031] = 141;
// bram[53032] = 165;
// bram[53033] = 187;
// bram[53034] = 208;
// bram[53035] = 225;
// bram[53036] = 238;
// bram[53037] = 248;
// bram[53038] = 253;
// bram[53039] = 253;
// bram[53040] = 248;
// bram[53041] = 239;
// bram[53042] = 226;
// bram[53043] = 209;
// bram[53044] = 189;
// bram[53045] = 166;
// bram[53046] = 143;
// bram[53047] = 118;
// bram[53048] = 94;
// bram[53049] = 71;
// bram[53050] = 50;
// bram[53051] = 32;
// bram[53052] = 17;
// bram[53053] = 7;
// bram[53054] = 1;
// bram[53055] = 0;
// bram[53056] = 3;
// bram[53057] = 11;
// bram[53058] = 24;
// bram[53059] = 40;
// bram[53060] = 59;
// bram[53061] = 81;
// bram[53062] = 105;
// bram[53063] = 129;
// bram[53064] = 154;
// bram[53065] = 177;
// bram[53066] = 199;
// bram[53067] = 217;
// bram[53068] = 233;
// bram[53069] = 244;
// bram[53070] = 251;
// bram[53071] = 253;
// bram[53072] = 251;
// bram[53073] = 244;
// bram[53074] = 233;
// bram[53075] = 217;
// bram[53076] = 198;
// bram[53077] = 177;
// bram[53078] = 154;
// bram[53079] = 129;
// bram[53080] = 105;
// bram[53081] = 81;
// bram[53082] = 59;
// bram[53083] = 40;
// bram[53084] = 23;
// bram[53085] = 11;
// bram[53086] = 3;
// bram[53087] = 0;
// bram[53088] = 1;
// bram[53089] = 7;
// bram[53090] = 17;
// bram[53091] = 32;
// bram[53092] = 50;
// bram[53093] = 71;
// bram[53094] = 94;
// bram[53095] = 118;
// bram[53096] = 143;
// bram[53097] = 167;
// bram[53098] = 189;
// bram[53099] = 209;
// bram[53100] = 226;
// bram[53101] = 239;
// bram[53102] = 249;
// bram[53103] = 253;
// bram[53104] = 253;
// bram[53105] = 248;
// bram[53106] = 238;
// bram[53107] = 225;
// bram[53108] = 207;
// bram[53109] = 187;
// bram[53110] = 164;
// bram[53111] = 140;
// bram[53112] = 116;
// bram[53113] = 92;
// bram[53114] = 69;
// bram[53115] = 48;
// bram[53116] = 30;
// bram[53117] = 16;
// bram[53118] = 6;
// bram[53119] = 1;
// bram[53120] = 0;
// bram[53121] = 4;
// bram[53122] = 12;
// bram[53123] = 25;
// bram[53124] = 41;
// bram[53125] = 61;
// bram[53126] = 83;
// bram[53127] = 107;
// bram[53128] = 132;
// bram[53129] = 156;
// bram[53130] = 179;
// bram[53131] = 200;
// bram[53132] = 219;
// bram[53133] = 234;
// bram[53134] = 245;
// bram[53135] = 252;
// bram[53136] = 253;
// bram[53137] = 251;
// bram[53138] = 243;
// bram[53139] = 231;
// bram[53140] = 216;
// bram[53141] = 197;
// bram[53142] = 175;
// bram[53143] = 151;
// bram[53144] = 127;
// bram[53145] = 102;
// bram[53146] = 79;
// bram[53147] = 57;
// bram[53148] = 38;
// bram[53149] = 22;
// bram[53150] = 10;
// bram[53151] = 3;
// bram[53152] = 0;
// bram[53153] = 1;
// bram[53154] = 8;
// bram[53155] = 19;
// bram[53156] = 34;
// bram[53157] = 52;
// bram[53158] = 73;
// bram[53159] = 96;
// bram[53160] = 121;
// bram[53161] = 145;
// bram[53162] = 169;
// bram[53163] = 191;
// bram[53164] = 211;
// bram[53165] = 228;
// bram[53166] = 241;
// bram[53167] = 249;
// bram[53168] = 253;
// bram[53169] = 253;
// bram[53170] = 247;
// bram[53171] = 237;
// bram[53172] = 223;
// bram[53173] = 206;
// bram[53174] = 185;
// bram[53175] = 162;
// bram[53176] = 138;
// bram[53177] = 114;
// bram[53178] = 89;
// bram[53179] = 67;
// bram[53180] = 46;
// bram[53181] = 29;
// bram[53182] = 15;
// bram[53183] = 5;
// bram[53184] = 0;
// bram[53185] = 0;
// bram[53186] = 4;
// bram[53187] = 13;
// bram[53188] = 26;
// bram[53189] = 43;
// bram[53190] = 63;
// bram[53191] = 86;
// bram[53192] = 109;
// bram[53193] = 134;
// bram[53194] = 158;
// bram[53195] = 181;
// bram[53196] = 202;
// bram[53197] = 220;
// bram[53198] = 235;
// bram[53199] = 246;
// bram[53200] = 252;
// bram[53201] = 253;
// bram[53202] = 250;
// bram[53203] = 242;
// bram[53204] = 230;
// bram[53205] = 214;
// bram[53206] = 195;
// bram[53207] = 173;
// bram[53208] = 149;
// bram[53209] = 125;
// bram[53210] = 100;
// bram[53211] = 77;
// bram[53212] = 55;
// bram[53213] = 36;
// bram[53214] = 21;
// bram[53215] = 9;
// bram[53216] = 2;
// bram[53217] = 0;
// bram[53218] = 2;
// bram[53219] = 9;
// bram[53220] = 20;
// bram[53221] = 35;
// bram[53222] = 54;
// bram[53223] = 75;
// bram[53224] = 98;
// bram[53225] = 123;
// bram[53226] = 147;
// bram[53227] = 171;
// bram[53228] = 193;
// bram[53229] = 213;
// bram[53230] = 229;
// bram[53231] = 241;
// bram[53232] = 250;
// bram[53233] = 253;
// bram[53234] = 252;
// bram[53235] = 246;
// bram[53236] = 236;
// bram[53237] = 222;
// bram[53238] = 204;
// bram[53239] = 183;
// bram[53240] = 160;
// bram[53241] = 136;
// bram[53242] = 111;
// bram[53243] = 87;
// bram[53244] = 65;
// bram[53245] = 45;
// bram[53246] = 27;
// bram[53247] = 14;
// bram[53248] = 5;
// bram[53249] = 0;
// bram[53250] = 0;
// bram[53251] = 5;
// bram[53252] = 14;
// bram[53253] = 28;
// bram[53254] = 45;
// bram[53255] = 65;
// bram[53256] = 88;
// bram[53257] = 112;
// bram[53258] = 136;
// bram[53259] = 160;
// bram[53260] = 183;
// bram[53261] = 204;
// bram[53262] = 222;
// bram[53263] = 236;
// bram[53264] = 247;
// bram[53265] = 252;
// bram[53266] = 253;
// bram[53267] = 250;
// bram[53268] = 241;
// bram[53269] = 229;
// bram[53270] = 212;
// bram[53271] = 193;
// bram[53272] = 171;
// bram[53273] = 147;
// bram[53274] = 122;
// bram[53275] = 98;
// bram[53276] = 75;
// bram[53277] = 53;
// bram[53278] = 35;
// bram[53279] = 20;
// bram[53280] = 8;
// bram[53281] = 2;
// bram[53282] = 0;
// bram[53283] = 2;
// bram[53284] = 9;
// bram[53285] = 21;
// bram[53286] = 37;
// bram[53287] = 56;
// bram[53288] = 77;
// bram[53289] = 101;
// bram[53290] = 125;
// bram[53291] = 149;
// bram[53292] = 173;
// bram[53293] = 195;
// bram[53294] = 214;
// bram[53295] = 230;
// bram[53296] = 242;
// bram[53297] = 250;
// bram[53298] = 253;
// bram[53299] = 252;
// bram[53300] = 246;
// bram[53301] = 235;
// bram[53302] = 220;
// bram[53303] = 202;
// bram[53304] = 181;
// bram[53305] = 158;
// bram[53306] = 134;
// bram[53307] = 109;
// bram[53308] = 85;
// bram[53309] = 63;
// bram[53310] = 43;
// bram[53311] = 26;
// bram[53312] = 13;
// bram[53313] = 4;
// bram[53314] = 0;
// bram[53315] = 0;
// bram[53316] = 6;
// bram[53317] = 15;
// bram[53318] = 29;
// bram[53319] = 47;
// bram[53320] = 67;
// bram[53321] = 90;
// bram[53322] = 114;
// bram[53323] = 138;
// bram[53324] = 163;
// bram[53325] = 185;
// bram[53326] = 206;
// bram[53327] = 223;
// bram[53328] = 237;
// bram[53329] = 247;
// bram[53330] = 253;
// bram[53331] = 253;
// bram[53332] = 249;
// bram[53333] = 240;
// bram[53334] = 227;
// bram[53335] = 211;
// bram[53336] = 191;
// bram[53337] = 169;
// bram[53338] = 145;
// bram[53339] = 120;
// bram[53340] = 96;
// bram[53341] = 73;
// bram[53342] = 52;
// bram[53343] = 33;
// bram[53344] = 18;
// bram[53345] = 8;
// bram[53346] = 1;
// bram[53347] = 0;
// bram[53348] = 3;
// bram[53349] = 10;
// bram[53350] = 22;
// bram[53351] = 38;
// bram[53352] = 57;
// bram[53353] = 79;
// bram[53354] = 103;
// bram[53355] = 127;
// bram[53356] = 152;
// bram[53357] = 175;
// bram[53358] = 197;
// bram[53359] = 216;
// bram[53360] = 232;
// bram[53361] = 243;
// bram[53362] = 251;
// bram[53363] = 253;
// bram[53364] = 252;
// bram[53365] = 245;
// bram[53366] = 234;
// bram[53367] = 219;
// bram[53368] = 200;
// bram[53369] = 179;
// bram[53370] = 156;
// bram[53371] = 131;
// bram[53372] = 107;
// bram[53373] = 83;
// bram[53374] = 61;
// bram[53375] = 41;
// bram[53376] = 25;
// bram[53377] = 12;
// bram[53378] = 4;
// bram[53379] = 0;
// bram[53380] = 1;
// bram[53381] = 6;
// bram[53382] = 16;
// bram[53383] = 31;
// bram[53384] = 48;
// bram[53385] = 69;
// bram[53386] = 92;
// bram[53387] = 116;
// bram[53388] = 141;
// bram[53389] = 165;
// bram[53390] = 187;
// bram[53391] = 208;
// bram[53392] = 225;
// bram[53393] = 238;
// bram[53394] = 248;
// bram[53395] = 253;
// bram[53396] = 253;
// bram[53397] = 248;
// bram[53398] = 239;
// bram[53399] = 226;
// bram[53400] = 209;
// bram[53401] = 189;
// bram[53402] = 166;
// bram[53403] = 142;
// bram[53404] = 118;
// bram[53405] = 94;
// bram[53406] = 71;
// bram[53407] = 50;
// bram[53408] = 32;
// bram[53409] = 17;
// bram[53410] = 7;
// bram[53411] = 1;
// bram[53412] = 0;
// bram[53413] = 3;
// bram[53414] = 11;
// bram[53415] = 24;
// bram[53416] = 40;
// bram[53417] = 59;
// bram[53418] = 81;
// bram[53419] = 105;
// bram[53420] = 129;
// bram[53421] = 154;
// bram[53422] = 177;
// bram[53423] = 199;
// bram[53424] = 217;
// bram[53425] = 233;
// bram[53426] = 244;
// bram[53427] = 251;
// bram[53428] = 253;
// bram[53429] = 251;
// bram[53430] = 244;
// bram[53431] = 233;
// bram[53432] = 217;
// bram[53433] = 198;
// bram[53434] = 177;
// bram[53435] = 153;
// bram[53436] = 129;
// bram[53437] = 105;
// bram[53438] = 81;
// bram[53439] = 59;
// bram[53440] = 40;
// bram[53441] = 23;
// bram[53442] = 11;
// bram[53443] = 3;
// bram[53444] = 0;
// bram[53445] = 1;
// bram[53446] = 7;
// bram[53447] = 17;
// bram[53448] = 32;
// bram[53449] = 50;
// bram[53450] = 71;
// bram[53451] = 94;
// bram[53452] = 118;
// bram[53453] = 143;
// bram[53454] = 167;
// bram[53455] = 189;
// bram[53456] = 209;
// bram[53457] = 226;
// bram[53458] = 240;
// bram[53459] = 249;
// bram[53460] = 253;
// bram[53461] = 253;
// bram[53462] = 248;
// bram[53463] = 238;
// bram[53464] = 225;
// bram[53465] = 207;
// bram[53466] = 187;
// bram[53467] = 164;
// bram[53468] = 140;
// bram[53469] = 116;
// bram[53470] = 92;
// bram[53471] = 69;
// bram[53472] = 48;
// bram[53473] = 30;
// bram[53474] = 16;
// bram[53475] = 6;
// bram[53476] = 1;
// bram[53477] = 0;
// bram[53478] = 4;
// bram[53479] = 12;
// bram[53480] = 25;
// bram[53481] = 42;
// bram[53482] = 61;
// bram[53483] = 83;
// bram[53484] = 107;
// bram[53485] = 132;
// bram[53486] = 156;
// bram[53487] = 179;
// bram[53488] = 201;
// bram[53489] = 219;
// bram[53490] = 234;
// bram[53491] = 245;
// bram[53492] = 252;
// bram[53493] = 253;
// bram[53494] = 251;
// bram[53495] = 243;
// bram[53496] = 231;
// bram[53497] = 216;
// bram[53498] = 196;
// bram[53499] = 175;
// bram[53500] = 151;
// bram[53501] = 127;
// bram[53502] = 102;
// bram[53503] = 79;
// bram[53504] = 57;
// bram[53505] = 38;
// bram[53506] = 22;
// bram[53507] = 10;
// bram[53508] = 3;
// bram[53509] = 0;
// bram[53510] = 1;
// bram[53511] = 8;
// bram[53512] = 19;
// bram[53513] = 34;
// bram[53514] = 52;
// bram[53515] = 73;
// bram[53516] = 96;
// bram[53517] = 121;
// bram[53518] = 145;
// bram[53519] = 169;
// bram[53520] = 191;
// bram[53521] = 211;
// bram[53522] = 228;
// bram[53523] = 241;
// bram[53524] = 249;
// bram[53525] = 253;
// bram[53526] = 253;
// bram[53527] = 247;
// bram[53528] = 237;
// bram[53529] = 223;
// bram[53530] = 206;
// bram[53531] = 185;
// bram[53532] = 162;
// bram[53533] = 138;
// bram[53534] = 113;
// bram[53535] = 89;
// bram[53536] = 67;
// bram[53537] = 46;
// bram[53538] = 29;
// bram[53539] = 15;
// bram[53540] = 5;
// bram[53541] = 0;
// bram[53542] = 0;
// bram[53543] = 4;
// bram[53544] = 13;
// bram[53545] = 26;
// bram[53546] = 43;
// bram[53547] = 63;
// bram[53548] = 86;
// bram[53549] = 109;
// bram[53550] = 134;
// bram[53551] = 158;
// bram[53552] = 181;
// bram[53553] = 202;
// bram[53554] = 221;
// bram[53555] = 235;
// bram[53556] = 246;
// bram[53557] = 252;
// bram[53558] = 253;
// bram[53559] = 250;
// bram[53560] = 242;
// bram[53561] = 230;
// bram[53562] = 214;
// bram[53563] = 195;
// bram[53564] = 173;
// bram[53565] = 149;
// bram[53566] = 125;
// bram[53567] = 100;
// bram[53568] = 77;
// bram[53569] = 55;
// bram[53570] = 36;
// bram[53571] = 21;
// bram[53572] = 9;
// bram[53573] = 2;
// bram[53574] = 0;
// bram[53575] = 2;
// bram[53576] = 9;
// bram[53577] = 20;
// bram[53578] = 35;
// bram[53579] = 54;
// bram[53580] = 75;
// bram[53581] = 98;
// bram[53582] = 123;
// bram[53583] = 147;
// bram[53584] = 171;
// bram[53585] = 193;
// bram[53586] = 213;
// bram[53587] = 229;
// bram[53588] = 241;
// bram[53589] = 250;
// bram[53590] = 253;
// bram[53591] = 252;
// bram[53592] = 246;
// bram[53593] = 236;
// bram[53594] = 222;
// bram[53595] = 204;
// bram[53596] = 183;
// bram[53597] = 160;
// bram[53598] = 136;
// bram[53599] = 111;
// bram[53600] = 87;
// bram[53601] = 65;
// bram[53602] = 45;
// bram[53603] = 27;
// bram[53604] = 14;
// bram[53605] = 5;
// bram[53606] = 0;
// bram[53607] = 0;
// bram[53608] = 5;
// bram[53609] = 14;
// bram[53610] = 28;
// bram[53611] = 45;
// bram[53612] = 65;
// bram[53613] = 88;
// bram[53614] = 112;
// bram[53615] = 136;
// bram[53616] = 160;
// bram[53617] = 183;
// bram[53618] = 204;
// bram[53619] = 222;
// bram[53620] = 236;
// bram[53621] = 247;
// bram[53622] = 252;
// bram[53623] = 253;
// bram[53624] = 250;
// bram[53625] = 241;
// bram[53626] = 229;
// bram[53627] = 212;
// bram[53628] = 193;
// bram[53629] = 171;
// bram[53630] = 147;
// bram[53631] = 122;
// bram[53632] = 98;
// bram[53633] = 75;
// bram[53634] = 53;
// bram[53635] = 35;
// bram[53636] = 20;
// bram[53637] = 8;
// bram[53638] = 2;
// bram[53639] = 0;
// bram[53640] = 2;
// bram[53641] = 9;
// bram[53642] = 21;
// bram[53643] = 37;
// bram[53644] = 56;
// bram[53645] = 77;
// bram[53646] = 101;
// bram[53647] = 125;
// bram[53648] = 150;
// bram[53649] = 173;
// bram[53650] = 195;
// bram[53651] = 214;
// bram[53652] = 230;
// bram[53653] = 242;
// bram[53654] = 250;
// bram[53655] = 253;
// bram[53656] = 252;
// bram[53657] = 246;
// bram[53658] = 235;
// bram[53659] = 220;
// bram[53660] = 202;
// bram[53661] = 181;
// bram[53662] = 158;
// bram[53663] = 134;
// bram[53664] = 109;
// bram[53665] = 85;
// bram[53666] = 63;
// bram[53667] = 43;
// bram[53668] = 26;
// bram[53669] = 13;
// bram[53670] = 4;
// bram[53671] = 0;
// bram[53672] = 0;
// bram[53673] = 6;
// bram[53674] = 15;
// bram[53675] = 29;
// bram[53676] = 47;
// bram[53677] = 67;
// bram[53678] = 90;
// bram[53679] = 114;
// bram[53680] = 138;
// bram[53681] = 163;
// bram[53682] = 185;
// bram[53683] = 206;
// bram[53684] = 223;
// bram[53685] = 237;
// bram[53686] = 247;
// bram[53687] = 253;
// bram[53688] = 253;
// bram[53689] = 249;
// bram[53690] = 240;
// bram[53691] = 227;
// bram[53692] = 211;
// bram[53693] = 191;
// bram[53694] = 168;
// bram[53695] = 145;
// bram[53696] = 120;
// bram[53697] = 96;
// bram[53698] = 73;
// bram[53699] = 52;
// bram[53700] = 33;
// bram[53701] = 18;
// bram[53702] = 8;
// bram[53703] = 1;
// bram[53704] = 0;
// bram[53705] = 3;
// bram[53706] = 10;
// bram[53707] = 22;
// bram[53708] = 38;
// bram[53709] = 57;
// bram[53710] = 79;
// bram[53711] = 103;
// bram[53712] = 127;
// bram[53713] = 152;
// bram[53714] = 175;
// bram[53715] = 197;
// bram[53716] = 216;
// bram[53717] = 232;
// bram[53718] = 243;
// bram[53719] = 251;
// bram[53720] = 253;
// bram[53721] = 251;
// bram[53722] = 245;
// bram[53723] = 234;
// bram[53724] = 219;
// bram[53725] = 200;
// bram[53726] = 179;
// bram[53727] = 156;
// bram[53728] = 131;
// bram[53729] = 107;
// bram[53730] = 83;
// bram[53731] = 61;
// bram[53732] = 41;
// bram[53733] = 25;
// bram[53734] = 12;
// bram[53735] = 4;
// bram[53736] = 0;
// bram[53737] = 1;
// bram[53738] = 6;
// bram[53739] = 16;
// bram[53740] = 31;
// bram[53741] = 48;
// bram[53742] = 69;
// bram[53743] = 92;
// bram[53744] = 116;
// bram[53745] = 141;
// bram[53746] = 165;
// bram[53747] = 187;
// bram[53748] = 208;
// bram[53749] = 225;
// bram[53750] = 239;
// bram[53751] = 248;
// bram[53752] = 253;
// bram[53753] = 253;
// bram[53754] = 248;
// bram[53755] = 239;
// bram[53756] = 226;
// bram[53757] = 209;
// bram[53758] = 189;
// bram[53759] = 166;
// bram[53760] = 142;
// bram[53761] = 118;
// bram[53762] = 94;
// bram[53763] = 71;
// bram[53764] = 50;
// bram[53765] = 32;
// bram[53766] = 17;
// bram[53767] = 7;
// bram[53768] = 1;
// bram[53769] = 0;
// bram[53770] = 3;
// bram[53771] = 11;
// bram[53772] = 24;
// bram[53773] = 40;
// bram[53774] = 59;
// bram[53775] = 81;
// bram[53776] = 105;
// bram[53777] = 130;
// bram[53778] = 154;
// bram[53779] = 177;
// bram[53780] = 199;
// bram[53781] = 217;
// bram[53782] = 233;
// bram[53783] = 244;
// bram[53784] = 251;
// bram[53785] = 253;
// bram[53786] = 251;
// bram[53787] = 244;
// bram[53788] = 233;
// bram[53789] = 217;
// bram[53790] = 198;
// bram[53791] = 177;
// bram[53792] = 153;
// bram[53793] = 129;
// bram[53794] = 105;
// bram[53795] = 81;
// bram[53796] = 59;
// bram[53797] = 40;
// bram[53798] = 23;
// bram[53799] = 11;
// bram[53800] = 3;
// bram[53801] = 0;
// bram[53802] = 1;
// bram[53803] = 7;
// bram[53804] = 17;
// bram[53805] = 32;
// bram[53806] = 50;
// bram[53807] = 71;
// bram[53808] = 94;
// bram[53809] = 118;
// bram[53810] = 143;
// bram[53811] = 167;
// bram[53812] = 189;
// bram[53813] = 209;
// bram[53814] = 226;
// bram[53815] = 240;
// bram[53816] = 249;
// bram[53817] = 253;
// bram[53818] = 253;
// bram[53819] = 248;
// bram[53820] = 238;
// bram[53821] = 225;
// bram[53822] = 207;
// bram[53823] = 187;
// bram[53824] = 164;
// bram[53825] = 140;
// bram[53826] = 116;
// bram[53827] = 91;
// bram[53828] = 69;
// bram[53829] = 48;
// bram[53830] = 30;
// bram[53831] = 16;
// bram[53832] = 6;
// bram[53833] = 1;
// bram[53834] = 0;
// bram[53835] = 4;
// bram[53836] = 12;
// bram[53837] = 25;
// bram[53838] = 42;
// bram[53839] = 61;
// bram[53840] = 83;
// bram[53841] = 107;
// bram[53842] = 132;
// bram[53843] = 156;
// bram[53844] = 179;
// bram[53845] = 201;
// bram[53846] = 219;
// bram[53847] = 234;
// bram[53848] = 245;
// bram[53849] = 252;
// bram[53850] = 253;
// bram[53851] = 251;
// bram[53852] = 243;
// bram[53853] = 231;
// bram[53854] = 216;
// bram[53855] = 196;
// bram[53856] = 175;
// bram[53857] = 151;
// bram[53858] = 127;
// bram[53859] = 102;
// bram[53860] = 79;
// bram[53861] = 57;
// bram[53862] = 38;
// bram[53863] = 22;
// bram[53864] = 10;
// bram[53865] = 3;
// bram[53866] = 0;
// bram[53867] = 1;
// bram[53868] = 8;
// bram[53869] = 19;
// bram[53870] = 34;
// bram[53871] = 52;
// bram[53872] = 73;
// bram[53873] = 96;
// bram[53874] = 121;
// bram[53875] = 145;
// bram[53876] = 169;
// bram[53877] = 191;
// bram[53878] = 211;
// bram[53879] = 228;
// bram[53880] = 241;
// bram[53881] = 249;
// bram[53882] = 253;
// bram[53883] = 253;
// bram[53884] = 247;
// bram[53885] = 237;
// bram[53886] = 223;
// bram[53887] = 205;
// bram[53888] = 185;
// bram[53889] = 162;
// bram[53890] = 138;
// bram[53891] = 113;
// bram[53892] = 89;
// bram[53893] = 67;
// bram[53894] = 46;
// bram[53895] = 29;
// bram[53896] = 15;
// bram[53897] = 5;
// bram[53898] = 0;
// bram[53899] = 0;
// bram[53900] = 4;
// bram[53901] = 13;
// bram[53902] = 26;
// bram[53903] = 43;
// bram[53904] = 63;
// bram[53905] = 86;
// bram[53906] = 109;
// bram[53907] = 134;
// bram[53908] = 158;
// bram[53909] = 181;
// bram[53910] = 202;
// bram[53911] = 221;
// bram[53912] = 235;
// bram[53913] = 246;
// bram[53914] = 252;
// bram[53915] = 253;
// bram[53916] = 250;
// bram[53917] = 242;
// bram[53918] = 230;
// bram[53919] = 214;
// bram[53920] = 195;
// bram[53921] = 173;
// bram[53922] = 149;
// bram[53923] = 125;
// bram[53924] = 100;
// bram[53925] = 77;
// bram[53926] = 55;
// bram[53927] = 36;
// bram[53928] = 21;
// bram[53929] = 9;
// bram[53930] = 2;
// bram[53931] = 0;
// bram[53932] = 2;
// bram[53933] = 9;
// bram[53934] = 20;
// bram[53935] = 35;
// bram[53936] = 54;
// bram[53937] = 75;
// bram[53938] = 99;
// bram[53939] = 123;
// bram[53940] = 147;
// bram[53941] = 171;
// bram[53942] = 193;
// bram[53943] = 213;
// bram[53944] = 229;
// bram[53945] = 242;
// bram[53946] = 250;
// bram[53947] = 253;
// bram[53948] = 252;
// bram[53949] = 246;
// bram[53950] = 236;
// bram[53951] = 222;
// bram[53952] = 204;
// bram[53953] = 183;
// bram[53954] = 160;
// bram[53955] = 136;
// bram[53956] = 111;
// bram[53957] = 87;
// bram[53958] = 65;
// bram[53959] = 45;
// bram[53960] = 27;
// bram[53961] = 14;
// bram[53962] = 5;
// bram[53963] = 0;
// bram[53964] = 0;
// bram[53965] = 5;
// bram[53966] = 14;
// bram[53967] = 28;
// bram[53968] = 45;
// bram[53969] = 65;
// bram[53970] = 88;
// bram[53971] = 112;
// bram[53972] = 136;
// bram[53973] = 160;
// bram[53974] = 183;
// bram[53975] = 204;
// bram[53976] = 222;
// bram[53977] = 236;
// bram[53978] = 247;
// bram[53979] = 252;
// bram[53980] = 253;
// bram[53981] = 250;
// bram[53982] = 241;
// bram[53983] = 229;
// bram[53984] = 212;
// bram[53985] = 193;
// bram[53986] = 171;
// bram[53987] = 147;
// bram[53988] = 122;
// bram[53989] = 98;
// bram[53990] = 75;
// bram[53991] = 53;
// bram[53992] = 35;
// bram[53993] = 20;
// bram[53994] = 8;
// bram[53995] = 2;
// bram[53996] = 0;
// bram[53997] = 2;
// bram[53998] = 9;
// bram[53999] = 21;
// bram[54000] = 37;
// bram[54001] = 56;
// bram[54002] = 77;
// bram[54003] = 101;
// bram[54004] = 125;
// bram[54005] = 150;
// bram[54006] = 173;
// bram[54007] = 195;
// bram[54008] = 214;
// bram[54009] = 230;
// bram[54010] = 242;
// bram[54011] = 250;
// bram[54012] = 253;
// bram[54013] = 252;
// bram[54014] = 246;
// bram[54015] = 235;
// bram[54016] = 220;
// bram[54017] = 202;
// bram[54018] = 181;
// bram[54019] = 158;
// bram[54020] = 133;
// bram[54021] = 109;
// bram[54022] = 85;
// bram[54023] = 63;
// bram[54024] = 43;
// bram[54025] = 26;
// bram[54026] = 13;
// bram[54027] = 4;
// bram[54028] = 0;
// bram[54029] = 0;
// bram[54030] = 6;
// bram[54031] = 15;
// bram[54032] = 29;
// bram[54033] = 47;
// bram[54034] = 67;
// bram[54035] = 90;
// bram[54036] = 114;
// bram[54037] = 139;
// bram[54038] = 163;
// bram[54039] = 185;
// bram[54040] = 206;
// bram[54041] = 223;
// bram[54042] = 237;
// bram[54043] = 247;
// bram[54044] = 253;
// bram[54045] = 253;
// bram[54046] = 249;
// bram[54047] = 240;
// bram[54048] = 227;
// bram[54049] = 211;
// bram[54050] = 191;
// bram[54051] = 168;
// bram[54052] = 145;
// bram[54053] = 120;
// bram[54054] = 96;
// bram[54055] = 73;
// bram[54056] = 52;
// bram[54057] = 33;
// bram[54058] = 18;
// bram[54059] = 8;
// bram[54060] = 1;
// bram[54061] = 0;
// bram[54062] = 3;
// bram[54063] = 10;
// bram[54064] = 22;
// bram[54065] = 38;
// bram[54066] = 58;
// bram[54067] = 79;
// bram[54068] = 103;
// bram[54069] = 127;
// bram[54070] = 152;
// bram[54071] = 175;
// bram[54072] = 197;
// bram[54073] = 216;
// bram[54074] = 232;
// bram[54075] = 243;
// bram[54076] = 251;
// bram[54077] = 253;
// bram[54078] = 251;
// bram[54079] = 245;
// bram[54080] = 234;
// bram[54081] = 219;
// bram[54082] = 200;
// bram[54083] = 179;
// bram[54084] = 156;
// bram[54085] = 131;
// bram[54086] = 107;
// bram[54087] = 83;
// bram[54088] = 61;
// bram[54089] = 41;
// bram[54090] = 25;
// bram[54091] = 12;
// bram[54092] = 4;
// bram[54093] = 0;
// bram[54094] = 1;
// bram[54095] = 6;
// bram[54096] = 16;
// bram[54097] = 31;
// bram[54098] = 48;
// bram[54099] = 69;
// bram[54100] = 92;
// bram[54101] = 116;
// bram[54102] = 141;
// bram[54103] = 165;
// bram[54104] = 187;
// bram[54105] = 208;
// bram[54106] = 225;
// bram[54107] = 239;
// bram[54108] = 248;
// bram[54109] = 253;
// bram[54110] = 253;
// bram[54111] = 248;
// bram[54112] = 239;
// bram[54113] = 226;
// bram[54114] = 209;
// bram[54115] = 189;
// bram[54116] = 166;
// bram[54117] = 142;
// bram[54118] = 118;
// bram[54119] = 94;
// bram[54120] = 71;
// bram[54121] = 50;
// bram[54122] = 32;
// bram[54123] = 17;
// bram[54124] = 7;
// bram[54125] = 1;
// bram[54126] = 0;
// bram[54127] = 3;
// bram[54128] = 11;
// bram[54129] = 24;
// bram[54130] = 40;
// bram[54131] = 59;
// bram[54132] = 81;
// bram[54133] = 105;
// bram[54134] = 130;
// bram[54135] = 154;
// bram[54136] = 177;
// bram[54137] = 199;
// bram[54138] = 217;
// bram[54139] = 233;
// bram[54140] = 244;
// bram[54141] = 251;
// bram[54142] = 253;
// bram[54143] = 251;
// bram[54144] = 244;
// bram[54145] = 233;
// bram[54146] = 217;
// bram[54147] = 198;
// bram[54148] = 177;
// bram[54149] = 153;
// bram[54150] = 129;
// bram[54151] = 105;
// bram[54152] = 81;
// bram[54153] = 59;
// bram[54154] = 39;
// bram[54155] = 23;
// bram[54156] = 11;
// bram[54157] = 3;
// bram[54158] = 0;
// bram[54159] = 1;
// bram[54160] = 7;
// bram[54161] = 18;
// bram[54162] = 32;
// bram[54163] = 50;
// bram[54164] = 71;
// bram[54165] = 94;
// bram[54166] = 118;
// bram[54167] = 143;
// bram[54168] = 167;
// bram[54169] = 189;
// bram[54170] = 209;
// bram[54171] = 226;
// bram[54172] = 240;
// bram[54173] = 249;
// bram[54174] = 253;
// bram[54175] = 253;
// bram[54176] = 248;
// bram[54177] = 238;
// bram[54178] = 225;
// bram[54179] = 207;
// bram[54180] = 187;
// bram[54181] = 164;
// bram[54182] = 140;
// bram[54183] = 116;
// bram[54184] = 91;
// bram[54185] = 69;
// bram[54186] = 48;
// bram[54187] = 30;
// bram[54188] = 16;
// bram[54189] = 6;
// bram[54190] = 1;
// bram[54191] = 0;
// bram[54192] = 4;
// bram[54193] = 12;
// bram[54194] = 25;
// bram[54195] = 42;
// bram[54196] = 61;
// bram[54197] = 84;
// bram[54198] = 107;
// bram[54199] = 132;
// bram[54200] = 156;
// bram[54201] = 179;
// bram[54202] = 201;
// bram[54203] = 219;
// bram[54204] = 234;
// bram[54205] = 245;
// bram[54206] = 252;
// bram[54207] = 253;
// bram[54208] = 251;
// bram[54209] = 243;
// bram[54210] = 231;
// bram[54211] = 215;
// bram[54212] = 196;
// bram[54213] = 175;
// bram[54214] = 151;
// bram[54215] = 127;
// bram[54216] = 102;
// bram[54217] = 79;
// bram[54218] = 57;
// bram[54219] = 38;
// bram[54220] = 22;
// bram[54221] = 10;
// bram[54222] = 2;
// bram[54223] = 0;
// bram[54224] = 1;
// bram[54225] = 8;
// bram[54226] = 19;
// bram[54227] = 34;
// bram[54228] = 52;
// bram[54229] = 73;
// bram[54230] = 96;
// bram[54231] = 121;
// bram[54232] = 145;
// bram[54233] = 169;
// bram[54234] = 191;
// bram[54235] = 211;
// bram[54236] = 228;
// bram[54237] = 241;
// bram[54238] = 249;
// bram[54239] = 253;
// bram[54240] = 252;
// bram[54241] = 247;
// bram[54242] = 237;
// bram[54243] = 223;
// bram[54244] = 205;
// bram[54245] = 185;
// bram[54246] = 162;
// bram[54247] = 138;
// bram[54248] = 113;
// bram[54249] = 89;
// bram[54250] = 67;
// bram[54251] = 46;
// bram[54252] = 29;
// bram[54253] = 15;
// bram[54254] = 5;
// bram[54255] = 0;
// bram[54256] = 0;
// bram[54257] = 4;
// bram[54258] = 13;
// bram[54259] = 26;
// bram[54260] = 43;
// bram[54261] = 63;
// bram[54262] = 86;
// bram[54263] = 110;
// bram[54264] = 134;
// bram[54265] = 158;
// bram[54266] = 181;
// bram[54267] = 202;
// bram[54268] = 221;
// bram[54269] = 235;
// bram[54270] = 246;
// bram[54271] = 252;
// bram[54272] = 253;
// bram[54273] = 250;
// bram[54274] = 242;
// bram[54275] = 230;
// bram[54276] = 214;
// bram[54277] = 195;
// bram[54278] = 173;
// bram[54279] = 149;
// bram[54280] = 125;
// bram[54281] = 100;
// bram[54282] = 77;
// bram[54283] = 55;
// bram[54284] = 36;
// bram[54285] = 21;
// bram[54286] = 9;
// bram[54287] = 2;
// bram[54288] = 0;
// bram[54289] = 2;
// bram[54290] = 9;
// bram[54291] = 20;
// bram[54292] = 35;
// bram[54293] = 54;
// bram[54294] = 75;
// bram[54295] = 99;
// bram[54296] = 123;
// bram[54297] = 147;
// bram[54298] = 171;
// bram[54299] = 193;
// bram[54300] = 213;
// bram[54301] = 229;
// bram[54302] = 242;
// bram[54303] = 250;
// bram[54304] = 253;
// bram[54305] = 252;
// bram[54306] = 246;
// bram[54307] = 236;
// bram[54308] = 222;
// bram[54309] = 204;
// bram[54310] = 183;
// bram[54311] = 160;
// bram[54312] = 136;
// bram[54313] = 111;
// bram[54314] = 87;
// bram[54315] = 65;
// bram[54316] = 44;
// bram[54317] = 27;
// bram[54318] = 14;
// bram[54319] = 5;
// bram[54320] = 0;
// bram[54321] = 0;
// bram[54322] = 5;
// bram[54323] = 14;
// bram[54324] = 28;
// bram[54325] = 45;
// bram[54326] = 65;
// bram[54327] = 88;
// bram[54328] = 112;
// bram[54329] = 136;
// bram[54330] = 160;
// bram[54331] = 183;
// bram[54332] = 204;
// bram[54333] = 222;
// bram[54334] = 236;
// bram[54335] = 247;
// bram[54336] = 252;
// bram[54337] = 253;
// bram[54338] = 250;
// bram[54339] = 241;
// bram[54340] = 229;
// bram[54341] = 212;
// bram[54342] = 193;
// bram[54343] = 171;
// bram[54344] = 147;
// bram[54345] = 122;
// bram[54346] = 98;
// bram[54347] = 75;
// bram[54348] = 53;
// bram[54349] = 35;
// bram[54350] = 20;
// bram[54351] = 8;
// bram[54352] = 2;
// bram[54353] = 0;
// bram[54354] = 2;
// bram[54355] = 9;
// bram[54356] = 21;
// bram[54357] = 37;
// bram[54358] = 56;
// bram[54359] = 77;
// bram[54360] = 101;
// bram[54361] = 125;
// bram[54362] = 150;
// bram[54363] = 173;
// bram[54364] = 195;
// bram[54365] = 214;
// bram[54366] = 230;
// bram[54367] = 242;
// bram[54368] = 250;
// bram[54369] = 253;
// bram[54370] = 252;
// bram[54371] = 246;
// bram[54372] = 235;
// bram[54373] = 220;
// bram[54374] = 202;
// bram[54375] = 181;
// bram[54376] = 158;
// bram[54377] = 133;
// bram[54378] = 109;
// bram[54379] = 85;
// bram[54380] = 63;
// bram[54381] = 43;
// bram[54382] = 26;
// bram[54383] = 13;
// bram[54384] = 4;
// bram[54385] = 0;
// bram[54386] = 0;
// bram[54387] = 6;
// bram[54388] = 15;
// bram[54389] = 29;
// bram[54390] = 47;
// bram[54391] = 67;
// bram[54392] = 90;
// bram[54393] = 114;
// bram[54394] = 139;
// bram[54395] = 163;
// bram[54396] = 185;
// bram[54397] = 206;
// bram[54398] = 224;
// bram[54399] = 237;
// bram[54400] = 247;
// bram[54401] = 253;
// bram[54402] = 253;
// bram[54403] = 249;
// bram[54404] = 240;
// bram[54405] = 227;
// bram[54406] = 211;
// bram[54407] = 191;
// bram[54408] = 168;
// bram[54409] = 145;
// bram[54410] = 120;
// bram[54411] = 96;
// bram[54412] = 73;
// bram[54413] = 51;
// bram[54414] = 33;
// bram[54415] = 18;
// bram[54416] = 8;
// bram[54417] = 1;
// bram[54418] = 0;
// bram[54419] = 3;
// bram[54420] = 10;
// bram[54421] = 22;
// bram[54422] = 38;
// bram[54423] = 58;
// bram[54424] = 79;
// bram[54425] = 103;
// bram[54426] = 127;
// bram[54427] = 152;
// bram[54428] = 175;
// bram[54429] = 197;
// bram[54430] = 216;
// bram[54431] = 232;
// bram[54432] = 243;
// bram[54433] = 251;
// bram[54434] = 253;
// bram[54435] = 251;
// bram[54436] = 245;
// bram[54437] = 234;
// bram[54438] = 219;
// bram[54439] = 200;
// bram[54440] = 179;
// bram[54441] = 156;
// bram[54442] = 131;
// bram[54443] = 107;
// bram[54444] = 83;
// bram[54445] = 61;
// bram[54446] = 41;
// bram[54447] = 25;
// bram[54448] = 12;
// bram[54449] = 4;
// bram[54450] = 0;
// bram[54451] = 1;
// bram[54452] = 6;
// bram[54453] = 16;
// bram[54454] = 31;
// bram[54455] = 48;
// bram[54456] = 69;
// bram[54457] = 92;
// bram[54458] = 116;
// bram[54459] = 141;
// bram[54460] = 165;
// bram[54461] = 187;
// bram[54462] = 208;
// bram[54463] = 225;
// bram[54464] = 239;
// bram[54465] = 248;
// bram[54466] = 253;
// bram[54467] = 253;
// bram[54468] = 248;
// bram[54469] = 239;
// bram[54470] = 226;
// bram[54471] = 209;
// bram[54472] = 189;
// bram[54473] = 166;
// bram[54474] = 142;
// bram[54475] = 118;
// bram[54476] = 94;
// bram[54477] = 71;
// bram[54478] = 50;
// bram[54479] = 32;
// bram[54480] = 17;
// bram[54481] = 7;
// bram[54482] = 1;
// bram[54483] = 0;
// bram[54484] = 3;
// bram[54485] = 11;
// bram[54486] = 24;
// bram[54487] = 40;
// bram[54488] = 59;
// bram[54489] = 81;
// bram[54490] = 105;
// bram[54491] = 130;
// bram[54492] = 154;
// bram[54493] = 177;
// bram[54494] = 199;
// bram[54495] = 218;
// bram[54496] = 233;
// bram[54497] = 244;
// bram[54498] = 251;
// bram[54499] = 253;
// bram[54500] = 251;
// bram[54501] = 244;
// bram[54502] = 232;
// bram[54503] = 217;
// bram[54504] = 198;
// bram[54505] = 177;
// bram[54506] = 153;
// bram[54507] = 129;
// bram[54508] = 104;
// bram[54509] = 81;
// bram[54510] = 59;
// bram[54511] = 39;
// bram[54512] = 23;
// bram[54513] = 11;
// bram[54514] = 3;
// bram[54515] = 0;
// bram[54516] = 1;
// bram[54517] = 7;
// bram[54518] = 18;
// bram[54519] = 32;
// bram[54520] = 50;
// bram[54521] = 71;
// bram[54522] = 94;
// bram[54523] = 118;
// bram[54524] = 143;
// bram[54525] = 167;
// bram[54526] = 189;
// bram[54527] = 209;
// bram[54528] = 226;
// bram[54529] = 240;
// bram[54530] = 249;
// bram[54531] = 253;
// bram[54532] = 253;
// bram[54533] = 248;
// bram[54534] = 238;
// bram[54535] = 225;
// bram[54536] = 207;
// bram[54537] = 187;
// bram[54538] = 164;
// bram[54539] = 140;
// bram[54540] = 116;
// bram[54541] = 91;
// bram[54542] = 69;
// bram[54543] = 48;
// bram[54544] = 30;
// bram[54545] = 16;
// bram[54546] = 6;
// bram[54547] = 1;
// bram[54548] = 0;
// bram[54549] = 4;
// bram[54550] = 12;
// bram[54551] = 25;
// bram[54552] = 42;
// bram[54553] = 61;
// bram[54554] = 84;
// bram[54555] = 107;
// bram[54556] = 132;
// bram[54557] = 156;
// bram[54558] = 179;
// bram[54559] = 201;
// bram[54560] = 219;
// bram[54561] = 234;
// bram[54562] = 245;
// bram[54563] = 252;
// bram[54564] = 253;
// bram[54565] = 251;
// bram[54566] = 243;
// bram[54567] = 231;
// bram[54568] = 215;
// bram[54569] = 196;
// bram[54570] = 175;
// bram[54571] = 151;
// bram[54572] = 127;
// bram[54573] = 102;
// bram[54574] = 79;
// bram[54575] = 57;
// bram[54576] = 38;
// bram[54577] = 22;
// bram[54578] = 10;
// bram[54579] = 2;
// bram[54580] = 0;
// bram[54581] = 1;
// bram[54582] = 8;
// bram[54583] = 19;
// bram[54584] = 34;
// bram[54585] = 52;
// bram[54586] = 73;
// bram[54587] = 96;
// bram[54588] = 121;
// bram[54589] = 145;
// bram[54590] = 169;
// bram[54591] = 191;
// bram[54592] = 211;
// bram[54593] = 228;
// bram[54594] = 241;
// bram[54595] = 249;
// bram[54596] = 253;
// bram[54597] = 252;
// bram[54598] = 247;
// bram[54599] = 237;
// bram[54600] = 223;
// bram[54601] = 205;
// bram[54602] = 185;
// bram[54603] = 162;
// bram[54604] = 138;
// bram[54605] = 113;
// bram[54606] = 89;
// bram[54607] = 67;
// bram[54608] = 46;
// bram[54609] = 29;
// bram[54610] = 15;
// bram[54611] = 5;
// bram[54612] = 0;
// bram[54613] = 0;
// bram[54614] = 4;
// bram[54615] = 13;
// bram[54616] = 26;
// bram[54617] = 43;
// bram[54618] = 63;
// bram[54619] = 86;
// bram[54620] = 110;
// bram[54621] = 134;
// bram[54622] = 158;
// bram[54623] = 181;
// bram[54624] = 202;
// bram[54625] = 221;
// bram[54626] = 235;
// bram[54627] = 246;
// bram[54628] = 252;
// bram[54629] = 253;
// bram[54630] = 250;
// bram[54631] = 242;
// bram[54632] = 230;
// bram[54633] = 214;
// bram[54634] = 194;
// bram[54635] = 173;
// bram[54636] = 149;
// bram[54637] = 124;
// bram[54638] = 100;
// bram[54639] = 77;
// bram[54640] = 55;
// bram[54641] = 36;
// bram[54642] = 21;
// bram[54643] = 9;
// bram[54644] = 2;
// bram[54645] = 0;
// bram[54646] = 2;
// bram[54647] = 9;
// bram[54648] = 20;
// bram[54649] = 35;
// bram[54650] = 54;
// bram[54651] = 75;
// bram[54652] = 99;
// bram[54653] = 123;
// bram[54654] = 147;
// bram[54655] = 171;
// bram[54656] = 193;
// bram[54657] = 213;
// bram[54658] = 229;
// bram[54659] = 242;
// bram[54660] = 250;
// bram[54661] = 253;
// bram[54662] = 252;
// bram[54663] = 246;
// bram[54664] = 236;
// bram[54665] = 222;
// bram[54666] = 204;
// bram[54667] = 183;
// bram[54668] = 160;
// bram[54669] = 136;
// bram[54670] = 111;
// bram[54671] = 87;
// bram[54672] = 65;
// bram[54673] = 44;
// bram[54674] = 27;
// bram[54675] = 14;
// bram[54676] = 5;
// bram[54677] = 0;
// bram[54678] = 0;
// bram[54679] = 5;
// bram[54680] = 14;
// bram[54681] = 28;
// bram[54682] = 45;
// bram[54683] = 65;
// bram[54684] = 88;
// bram[54685] = 112;
// bram[54686] = 136;
// bram[54687] = 161;
// bram[54688] = 183;
// bram[54689] = 204;
// bram[54690] = 222;
// bram[54691] = 236;
// bram[54692] = 247;
// bram[54693] = 252;
// bram[54694] = 253;
// bram[54695] = 250;
// bram[54696] = 241;
// bram[54697] = 229;
// bram[54698] = 212;
// bram[54699] = 193;
// bram[54700] = 170;
// bram[54701] = 147;
// bram[54702] = 122;
// bram[54703] = 98;
// bram[54704] = 75;
// bram[54705] = 53;
// bram[54706] = 35;
// bram[54707] = 20;
// bram[54708] = 8;
// bram[54709] = 2;
// bram[54710] = 0;
// bram[54711] = 2;
// bram[54712] = 9;
// bram[54713] = 21;
// bram[54714] = 37;
// bram[54715] = 56;
// bram[54716] = 77;
// bram[54717] = 101;
// bram[54718] = 125;
// bram[54719] = 150;
// bram[54720] = 173;
// bram[54721] = 195;
// bram[54722] = 214;
// bram[54723] = 230;
// bram[54724] = 242;
// bram[54725] = 250;
// bram[54726] = 253;
// bram[54727] = 252;
// bram[54728] = 246;
// bram[54729] = 235;
// bram[54730] = 220;
// bram[54731] = 202;
// bram[54732] = 181;
// bram[54733] = 158;
// bram[54734] = 133;
// bram[54735] = 109;
// bram[54736] = 85;
// bram[54737] = 63;
// bram[54738] = 43;
// bram[54739] = 26;
// bram[54740] = 13;
// bram[54741] = 4;
// bram[54742] = 0;
// bram[54743] = 0;
// bram[54744] = 6;
// bram[54745] = 15;
// bram[54746] = 29;
// bram[54747] = 47;
// bram[54748] = 67;
// bram[54749] = 90;
// bram[54750] = 114;
// bram[54751] = 139;
// bram[54752] = 163;
// bram[54753] = 185;
// bram[54754] = 206;
// bram[54755] = 224;
// bram[54756] = 238;
// bram[54757] = 247;
// bram[54758] = 253;
// bram[54759] = 253;
// bram[54760] = 249;
// bram[54761] = 240;
// bram[54762] = 227;
// bram[54763] = 211;
// bram[54764] = 191;
// bram[54765] = 168;
// bram[54766] = 144;
// bram[54767] = 120;
// bram[54768] = 96;
// bram[54769] = 73;
// bram[54770] = 51;
// bram[54771] = 33;
// bram[54772] = 18;
// bram[54773] = 8;
// bram[54774] = 1;
// bram[54775] = 0;
// bram[54776] = 3;
// bram[54777] = 10;
// bram[54778] = 22;
// bram[54779] = 38;
// bram[54780] = 58;
// bram[54781] = 79;
// bram[54782] = 103;
// bram[54783] = 127;
// bram[54784] = 152;
// bram[54785] = 175;
// bram[54786] = 197;
// bram[54787] = 216;
// bram[54788] = 232;
// bram[54789] = 243;
// bram[54790] = 251;
// bram[54791] = 253;
// bram[54792] = 251;
// bram[54793] = 245;
// bram[54794] = 234;
// bram[54795] = 219;
// bram[54796] = 200;
// bram[54797] = 179;
// bram[54798] = 155;
// bram[54799] = 131;
// bram[54800] = 107;
// bram[54801] = 83;
// bram[54802] = 61;
// bram[54803] = 41;
// bram[54804] = 25;
// bram[54805] = 12;
// bram[54806] = 4;
// bram[54807] = 0;
// bram[54808] = 1;
// bram[54809] = 6;
// bram[54810] = 16;
// bram[54811] = 31;
// bram[54812] = 49;
// bram[54813] = 69;
// bram[54814] = 92;
// bram[54815] = 116;
// bram[54816] = 141;
// bram[54817] = 165;
// bram[54818] = 187;
// bram[54819] = 208;
// bram[54820] = 225;
// bram[54821] = 239;
// bram[54822] = 248;
// bram[54823] = 253;
// bram[54824] = 253;
// bram[54825] = 248;
// bram[54826] = 239;
// bram[54827] = 226;
// bram[54828] = 209;
// bram[54829] = 189;
// bram[54830] = 166;
// bram[54831] = 142;
// bram[54832] = 118;
// bram[54833] = 94;
// bram[54834] = 71;
// bram[54835] = 50;
// bram[54836] = 32;
// bram[54837] = 17;
// bram[54838] = 7;
// bram[54839] = 1;
// bram[54840] = 0;
// bram[54841] = 3;
// bram[54842] = 11;
// bram[54843] = 24;
// bram[54844] = 40;
// bram[54845] = 60;
// bram[54846] = 82;
// bram[54847] = 105;
// bram[54848] = 130;
// bram[54849] = 154;
// bram[54850] = 177;
// bram[54851] = 199;
// bram[54852] = 218;
// bram[54853] = 233;
// bram[54854] = 244;
// bram[54855] = 251;
// bram[54856] = 253;
// bram[54857] = 251;
// bram[54858] = 244;
// bram[54859] = 232;
// bram[54860] = 217;
// bram[54861] = 198;
// bram[54862] = 177;
// bram[54863] = 153;
// bram[54864] = 129;
// bram[54865] = 104;
// bram[54866] = 81;
// bram[54867] = 59;
// bram[54868] = 39;
// bram[54869] = 23;
// bram[54870] = 11;
// bram[54871] = 3;
// bram[54872] = 0;
// bram[54873] = 1;
// bram[54874] = 7;
// bram[54875] = 18;
// bram[54876] = 32;
// bram[54877] = 50;
// bram[54878] = 71;
// bram[54879] = 94;
// bram[54880] = 119;
// bram[54881] = 143;
// bram[54882] = 167;
// bram[54883] = 189;
// bram[54884] = 209;
// bram[54885] = 226;
// bram[54886] = 240;
// bram[54887] = 249;
// bram[54888] = 253;
// bram[54889] = 253;
// bram[54890] = 248;
// bram[54891] = 238;
// bram[54892] = 224;
// bram[54893] = 207;
// bram[54894] = 187;
// bram[54895] = 164;
// bram[54896] = 140;
// bram[54897] = 115;
// bram[54898] = 91;
// bram[54899] = 69;
// bram[54900] = 48;
// bram[54901] = 30;
// bram[54902] = 16;
// bram[54903] = 6;
// bram[54904] = 1;
// bram[54905] = 0;
// bram[54906] = 4;
// bram[54907] = 12;
// bram[54908] = 25;
// bram[54909] = 42;
// bram[54910] = 61;
// bram[54911] = 84;
// bram[54912] = 107;
// bram[54913] = 132;
// bram[54914] = 156;
// bram[54915] = 179;
// bram[54916] = 201;
// bram[54917] = 219;
// bram[54918] = 234;
// bram[54919] = 245;
// bram[54920] = 252;
// bram[54921] = 253;
// bram[54922] = 251;
// bram[54923] = 243;
// bram[54924] = 231;
// bram[54925] = 215;
// bram[54926] = 196;
// bram[54927] = 175;
// bram[54928] = 151;
// bram[54929] = 127;
// bram[54930] = 102;
// bram[54931] = 79;
// bram[54932] = 57;
// bram[54933] = 38;
// bram[54934] = 22;
// bram[54935] = 10;
// bram[54936] = 2;
// bram[54937] = 0;
// bram[54938] = 1;
// bram[54939] = 8;
// bram[54940] = 19;
// bram[54941] = 34;
// bram[54942] = 52;
// bram[54943] = 73;
// bram[54944] = 96;
// bram[54945] = 121;
// bram[54946] = 145;
// bram[54947] = 169;
// bram[54948] = 191;
// bram[54949] = 211;
// bram[54950] = 228;
// bram[54951] = 241;
// bram[54952] = 249;
// bram[54953] = 253;
// bram[54954] = 252;
// bram[54955] = 247;
// bram[54956] = 237;
// bram[54957] = 223;
// bram[54958] = 205;
// bram[54959] = 185;
// bram[54960] = 162;
// bram[54961] = 138;
// bram[54962] = 113;
// bram[54963] = 89;
// bram[54964] = 67;
// bram[54965] = 46;
// bram[54966] = 29;
// bram[54967] = 15;
// bram[54968] = 5;
// bram[54969] = 0;
// bram[54970] = 0;
// bram[54971] = 4;
// bram[54972] = 13;
// bram[54973] = 26;
// bram[54974] = 43;
// bram[54975] = 63;
// bram[54976] = 86;
// bram[54977] = 110;
// bram[54978] = 134;
// bram[54979] = 158;
// bram[54980] = 181;
// bram[54981] = 202;
// bram[54982] = 221;
// bram[54983] = 235;
// bram[54984] = 246;
// bram[54985] = 252;
// bram[54986] = 253;
// bram[54987] = 250;
// bram[54988] = 242;
// bram[54989] = 230;
// bram[54990] = 214;
// bram[54991] = 194;
// bram[54992] = 173;
// bram[54993] = 149;
// bram[54994] = 124;
// bram[54995] = 100;
// bram[54996] = 77;
// bram[54997] = 55;
// bram[54998] = 36;
// bram[54999] = 21;
// bram[55000] = 9;
// bram[55001] = 2;
// bram[55002] = 0;
// bram[55003] = 2;
// bram[55004] = 9;
// bram[55005] = 20;
// bram[55006] = 35;
// bram[55007] = 54;
// bram[55008] = 75;
// bram[55009] = 99;
// bram[55010] = 123;
// bram[55011] = 147;
// bram[55012] = 171;
// bram[55013] = 193;
// bram[55014] = 213;
// bram[55015] = 229;
// bram[55016] = 242;
// bram[55017] = 250;
// bram[55018] = 253;
// bram[55019] = 252;
// bram[55020] = 246;
// bram[55021] = 236;
// bram[55022] = 222;
// bram[55023] = 204;
// bram[55024] = 183;
// bram[55025] = 160;
// bram[55026] = 136;
// bram[55027] = 111;
// bram[55028] = 87;
// bram[55029] = 65;
// bram[55030] = 44;
// bram[55031] = 27;
// bram[55032] = 14;
// bram[55033] = 5;
// bram[55034] = 0;
// bram[55035] = 0;
// bram[55036] = 5;
// bram[55037] = 14;
// bram[55038] = 28;
// bram[55039] = 45;
// bram[55040] = 65;
// bram[55041] = 88;
// bram[55042] = 112;
// bram[55043] = 136;
// bram[55044] = 161;
// bram[55045] = 183;
// bram[55046] = 204;
// bram[55047] = 222;
// bram[55048] = 236;
// bram[55049] = 247;
// bram[55050] = 252;
// bram[55051] = 253;
// bram[55052] = 250;
// bram[55053] = 241;
// bram[55054] = 229;
// bram[55055] = 212;
// bram[55056] = 193;
// bram[55057] = 170;
// bram[55058] = 147;
// bram[55059] = 122;
// bram[55060] = 98;
// bram[55061] = 75;
// bram[55062] = 53;
// bram[55063] = 35;
// bram[55064] = 19;
// bram[55065] = 8;
// bram[55066] = 2;
// bram[55067] = 0;
// bram[55068] = 2;
// bram[55069] = 9;
// bram[55070] = 21;
// bram[55071] = 37;
// bram[55072] = 56;
// bram[55073] = 77;
// bram[55074] = 101;
// bram[55075] = 125;
// bram[55076] = 150;
// bram[55077] = 173;
// bram[55078] = 195;
// bram[55079] = 214;
// bram[55080] = 230;
// bram[55081] = 243;
// bram[55082] = 250;
// bram[55083] = 253;
// bram[55084] = 252;
// bram[55085] = 246;
// bram[55086] = 235;
// bram[55087] = 220;
// bram[55088] = 202;
// bram[55089] = 181;
// bram[55090] = 158;
// bram[55091] = 133;
// bram[55092] = 109;
// bram[55093] = 85;
// bram[55094] = 63;
// bram[55095] = 43;
// bram[55096] = 26;
// bram[55097] = 13;
// bram[55098] = 4;
// bram[55099] = 0;
// bram[55100] = 0;
// bram[55101] = 6;
// bram[55102] = 15;
// bram[55103] = 29;
// bram[55104] = 47;
// bram[55105] = 67;
// bram[55106] = 90;
// bram[55107] = 114;
// bram[55108] = 139;
// bram[55109] = 163;
// bram[55110] = 185;
// bram[55111] = 206;
// bram[55112] = 224;
// bram[55113] = 238;
// bram[55114] = 247;
// bram[55115] = 253;
// bram[55116] = 253;
// bram[55117] = 249;
// bram[55118] = 240;
// bram[55119] = 227;
// bram[55120] = 210;
// bram[55121] = 191;
// bram[55122] = 168;
// bram[55123] = 144;
// bram[55124] = 120;
// bram[55125] = 96;
// bram[55126] = 73;
// bram[55127] = 51;
// bram[55128] = 33;
// bram[55129] = 18;
// bram[55130] = 8;
// bram[55131] = 1;
// bram[55132] = 0;
// bram[55133] = 3;
// bram[55134] = 10;
// bram[55135] = 22;
// bram[55136] = 38;
// bram[55137] = 58;
// bram[55138] = 79;
// bram[55139] = 103;
// bram[55140] = 127;
// bram[55141] = 152;
// bram[55142] = 175;
// bram[55143] = 197;
// bram[55144] = 216;
// bram[55145] = 232;
// bram[55146] = 243;
// bram[55147] = 251;
// bram[55148] = 253;
// bram[55149] = 251;
// bram[55150] = 245;
// bram[55151] = 234;
// bram[55152] = 219;
// bram[55153] = 200;
// bram[55154] = 179;
// bram[55155] = 155;
// bram[55156] = 131;
// bram[55157] = 107;
// bram[55158] = 83;
// bram[55159] = 61;
// bram[55160] = 41;
// bram[55161] = 25;
// bram[55162] = 12;
// bram[55163] = 4;
// bram[55164] = 0;
// bram[55165] = 1;
// bram[55166] = 6;
// bram[55167] = 16;
// bram[55168] = 31;
// bram[55169] = 49;
// bram[55170] = 69;
// bram[55171] = 92;
// bram[55172] = 116;
// bram[55173] = 141;
// bram[55174] = 165;
// bram[55175] = 187;
// bram[55176] = 208;
// bram[55177] = 225;
// bram[55178] = 239;
// bram[55179] = 248;
// bram[55180] = 253;
// bram[55181] = 253;
// bram[55182] = 248;
// bram[55183] = 239;
// bram[55184] = 226;
// bram[55185] = 209;
// bram[55186] = 189;
// bram[55187] = 166;
// bram[55188] = 142;
// bram[55189] = 118;
// bram[55190] = 93;
// bram[55191] = 70;
// bram[55192] = 50;
// bram[55193] = 32;
// bram[55194] = 17;
// bram[55195] = 7;
// bram[55196] = 1;
// bram[55197] = 0;
// bram[55198] = 3;
// bram[55199] = 11;
// bram[55200] = 24;
// bram[55201] = 40;
// bram[55202] = 60;
// bram[55203] = 82;
// bram[55204] = 105;
// bram[55205] = 130;
// bram[55206] = 154;
// bram[55207] = 177;
// bram[55208] = 199;
// bram[55209] = 218;
// bram[55210] = 233;
// bram[55211] = 244;
// bram[55212] = 251;
// bram[55213] = 253;
// bram[55214] = 251;
// bram[55215] = 244;
// bram[55216] = 232;
// bram[55217] = 217;
// bram[55218] = 198;
// bram[55219] = 177;
// bram[55220] = 153;
// bram[55221] = 129;
// bram[55222] = 104;
// bram[55223] = 81;
// bram[55224] = 59;
// bram[55225] = 39;
// bram[55226] = 23;
// bram[55227] = 11;
// bram[55228] = 3;
// bram[55229] = 0;
// bram[55230] = 1;
// bram[55231] = 7;
// bram[55232] = 18;
// bram[55233] = 32;
// bram[55234] = 50;
// bram[55235] = 71;
// bram[55236] = 94;
// bram[55237] = 119;
// bram[55238] = 143;
// bram[55239] = 167;
// bram[55240] = 189;
// bram[55241] = 209;
// bram[55242] = 226;
// bram[55243] = 240;
// bram[55244] = 249;
// bram[55245] = 253;
// bram[55246] = 253;
// bram[55247] = 248;
// bram[55248] = 238;
// bram[55249] = 224;
// bram[55250] = 207;
// bram[55251] = 187;
// bram[55252] = 164;
// bram[55253] = 140;
// bram[55254] = 115;
// bram[55255] = 91;
// bram[55256] = 68;
// bram[55257] = 48;
// bram[55258] = 30;
// bram[55259] = 16;
// bram[55260] = 6;
// bram[55261] = 1;
// bram[55262] = 0;
// bram[55263] = 4;
// bram[55264] = 12;
// bram[55265] = 25;
// bram[55266] = 42;
// bram[55267] = 61;
// bram[55268] = 84;
// bram[55269] = 107;
// bram[55270] = 132;
// bram[55271] = 156;
// bram[55272] = 179;
// bram[55273] = 201;
// bram[55274] = 219;
// bram[55275] = 234;
// bram[55276] = 245;
// bram[55277] = 252;
// bram[55278] = 253;
// bram[55279] = 251;
// bram[55280] = 243;
// bram[55281] = 231;
// bram[55282] = 215;
// bram[55283] = 196;
// bram[55284] = 175;
// bram[55285] = 151;
// bram[55286] = 127;
// bram[55287] = 102;
// bram[55288] = 79;
// bram[55289] = 57;
// bram[55290] = 38;
// bram[55291] = 22;
// bram[55292] = 10;
// bram[55293] = 2;
// bram[55294] = 0;
// bram[55295] = 1;
// bram[55296] = 8;
// bram[55297] = 19;
// bram[55298] = 34;
// bram[55299] = 52;
// bram[55300] = 73;
// bram[55301] = 97;
// bram[55302] = 121;
// bram[55303] = 145;
// bram[55304] = 169;
// bram[55305] = 191;
// bram[55306] = 211;
// bram[55307] = 228;
// bram[55308] = 241;
// bram[55309] = 249;
// bram[55310] = 253;
// bram[55311] = 252;
// bram[55312] = 247;
// bram[55313] = 237;
// bram[55314] = 223;
// bram[55315] = 205;
// bram[55316] = 185;
// bram[55317] = 162;
// bram[55318] = 138;
// bram[55319] = 113;
// bram[55320] = 89;
// bram[55321] = 67;
// bram[55322] = 46;
// bram[55323] = 29;
// bram[55324] = 15;
// bram[55325] = 5;
// bram[55326] = 0;
// bram[55327] = 0;
// bram[55328] = 4;
// bram[55329] = 13;
// bram[55330] = 26;
// bram[55331] = 43;
// bram[55332] = 63;
// bram[55333] = 86;
// bram[55334] = 110;
// bram[55335] = 134;
// bram[55336] = 158;
// bram[55337] = 182;
// bram[55338] = 203;
// bram[55339] = 221;
// bram[55340] = 235;
// bram[55341] = 246;
// bram[55342] = 252;
// bram[55343] = 253;
// bram[55344] = 250;
// bram[55345] = 242;
// bram[55346] = 230;
// bram[55347] = 214;
// bram[55348] = 194;
// bram[55349] = 172;
// bram[55350] = 149;
// bram[55351] = 124;
// bram[55352] = 100;
// bram[55353] = 77;
// bram[55354] = 55;
// bram[55355] = 36;
// bram[55356] = 21;
// bram[55357] = 9;
// bram[55358] = 2;
// bram[55359] = 0;
// bram[55360] = 2;
// bram[55361] = 9;
// bram[55362] = 20;
// bram[55363] = 35;
// bram[55364] = 54;
// bram[55365] = 75;
// bram[55366] = 99;
// bram[55367] = 123;
// bram[55368] = 148;
// bram[55369] = 171;
// bram[55370] = 193;
// bram[55371] = 213;
// bram[55372] = 229;
// bram[55373] = 242;
// bram[55374] = 250;
// bram[55375] = 253;
// bram[55376] = 252;
// bram[55377] = 246;
// bram[55378] = 236;
// bram[55379] = 222;
// bram[55380] = 204;
// bram[55381] = 183;
// bram[55382] = 160;
// bram[55383] = 136;
// bram[55384] = 111;
// bram[55385] = 87;
// bram[55386] = 65;
// bram[55387] = 44;
// bram[55388] = 27;
// bram[55389] = 14;
// bram[55390] = 5;
// bram[55391] = 0;
// bram[55392] = 0;
// bram[55393] = 5;
// bram[55394] = 14;
// bram[55395] = 28;
// bram[55396] = 45;
// bram[55397] = 65;
// bram[55398] = 88;
// bram[55399] = 112;
// bram[55400] = 136;
// bram[55401] = 161;
// bram[55402] = 184;
// bram[55403] = 204;
// bram[55404] = 222;
// bram[55405] = 236;
// bram[55406] = 247;
// bram[55407] = 252;
// bram[55408] = 253;
// bram[55409] = 250;
// bram[55410] = 241;
// bram[55411] = 229;
// bram[55412] = 212;
// bram[55413] = 192;
// bram[55414] = 170;
// bram[55415] = 147;
// bram[55416] = 122;
// bram[55417] = 98;
// bram[55418] = 75;
// bram[55419] = 53;
// bram[55420] = 35;
// bram[55421] = 19;
// bram[55422] = 8;
// bram[55423] = 2;
// bram[55424] = 0;
// bram[55425] = 2;
// bram[55426] = 10;
// bram[55427] = 21;
// bram[55428] = 37;
// bram[55429] = 56;
// bram[55430] = 77;
// bram[55431] = 101;
// bram[55432] = 125;
// bram[55433] = 150;
// bram[55434] = 173;
// bram[55435] = 195;
// bram[55436] = 214;
// bram[55437] = 230;
// bram[55438] = 243;
// bram[55439] = 250;
// bram[55440] = 253;
// bram[55441] = 252;
// bram[55442] = 246;
// bram[55443] = 235;
// bram[55444] = 220;
// bram[55445] = 202;
// bram[55446] = 181;
// bram[55447] = 158;
// bram[55448] = 133;
// bram[55449] = 109;
// bram[55450] = 85;
// bram[55451] = 63;
// bram[55452] = 43;
// bram[55453] = 26;
// bram[55454] = 13;
// bram[55455] = 4;
// bram[55456] = 0;
// bram[55457] = 0;
// bram[55458] = 6;
// bram[55459] = 15;
// bram[55460] = 29;
// bram[55461] = 47;
// bram[55462] = 67;
// bram[55463] = 90;
// bram[55464] = 114;
// bram[55465] = 139;
// bram[55466] = 163;
// bram[55467] = 186;
// bram[55468] = 206;
// bram[55469] = 224;
// bram[55470] = 238;
// bram[55471] = 247;
// bram[55472] = 253;
// bram[55473] = 253;
// bram[55474] = 249;
// bram[55475] = 240;
// bram[55476] = 227;
// bram[55477] = 210;
// bram[55478] = 191;
// bram[55479] = 168;
// bram[55480] = 144;
// bram[55481] = 120;
// bram[55482] = 96;
// bram[55483] = 72;
// bram[55484] = 51;
// bram[55485] = 33;
// bram[55486] = 18;
// bram[55487] = 8;
// bram[55488] = 1;
// bram[55489] = 0;
// bram[55490] = 3;
// bram[55491] = 10;
// bram[55492] = 22;
// bram[55493] = 38;
// bram[55494] = 58;
// bram[55495] = 80;
// bram[55496] = 103;
// bram[55497] = 128;
// bram[55498] = 152;
// bram[55499] = 175;
// bram[55500] = 197;
// bram[55501] = 216;
// bram[55502] = 232;
// bram[55503] = 243;
// bram[55504] = 251;
// bram[55505] = 253;
// bram[55506] = 251;
// bram[55507] = 245;
// bram[55508] = 234;
// bram[55509] = 218;
// bram[55510] = 200;
// bram[55511] = 179;
// bram[55512] = 155;
// bram[55513] = 131;
// bram[55514] = 107;
// bram[55515] = 83;
// bram[55516] = 61;
// bram[55517] = 41;
// bram[55518] = 25;
// bram[55519] = 12;
// bram[55520] = 3;
// bram[55521] = 0;
// bram[55522] = 1;
// bram[55523] = 6;
// bram[55524] = 16;
// bram[55525] = 31;
// bram[55526] = 49;
// bram[55527] = 69;
// bram[55528] = 92;
// bram[55529] = 116;
// bram[55530] = 141;
// bram[55531] = 165;
// bram[55532] = 188;
// bram[55533] = 208;
// bram[55534] = 225;
// bram[55535] = 239;
// bram[55536] = 248;
// bram[55537] = 253;
// bram[55538] = 253;
// bram[55539] = 248;
// bram[55540] = 239;
// bram[55541] = 226;
// bram[55542] = 209;
// bram[55543] = 189;
// bram[55544] = 166;
// bram[55545] = 142;
// bram[55546] = 118;
// bram[55547] = 93;
// bram[55548] = 70;
// bram[55549] = 50;
// bram[55550] = 32;
// bram[55551] = 17;
// bram[55552] = 7;
// bram[55553] = 1;
// bram[55554] = 0;
// bram[55555] = 3;
// bram[55556] = 11;
// bram[55557] = 24;
// bram[55558] = 40;
// bram[55559] = 60;
// bram[55560] = 82;
// bram[55561] = 105;
// bram[55562] = 130;
// bram[55563] = 154;
// bram[55564] = 177;
// bram[55565] = 199;
// bram[55566] = 218;
// bram[55567] = 233;
// bram[55568] = 244;
// bram[55569] = 251;
// bram[55570] = 253;
// bram[55571] = 251;
// bram[55572] = 244;
// bram[55573] = 232;
// bram[55574] = 217;
// bram[55575] = 198;
// bram[55576] = 177;
// bram[55577] = 153;
// bram[55578] = 129;
// bram[55579] = 104;
// bram[55580] = 81;
// bram[55581] = 59;
// bram[55582] = 39;
// bram[55583] = 23;
// bram[55584] = 11;
// bram[55585] = 3;
// bram[55586] = 0;
// bram[55587] = 1;
// bram[55588] = 7;
// bram[55589] = 18;
// bram[55590] = 32;
// bram[55591] = 50;
// bram[55592] = 71;
// bram[55593] = 94;
// bram[55594] = 119;
// bram[55595] = 143;
// bram[55596] = 167;
// bram[55597] = 189;
// bram[55598] = 210;
// bram[55599] = 226;
// bram[55600] = 240;
// bram[55601] = 249;
// bram[55602] = 253;
// bram[55603] = 253;
// bram[55604] = 248;
// bram[55605] = 238;
// bram[55606] = 224;
// bram[55607] = 207;
// bram[55608] = 187;
// bram[55609] = 164;
// bram[55610] = 140;
// bram[55611] = 115;
// bram[55612] = 91;
// bram[55613] = 68;
// bram[55614] = 48;
// bram[55615] = 30;
// bram[55616] = 16;
// bram[55617] = 6;
// bram[55618] = 1;
// bram[55619] = 0;
// bram[55620] = 4;
// bram[55621] = 12;
// bram[55622] = 25;
// bram[55623] = 42;
// bram[55624] = 62;
// bram[55625] = 84;
// bram[55626] = 108;
// bram[55627] = 132;
// bram[55628] = 156;
// bram[55629] = 180;
// bram[55630] = 201;
// bram[55631] = 219;
// bram[55632] = 234;
// bram[55633] = 245;
// bram[55634] = 252;
// bram[55635] = 253;
// bram[55636] = 251;
// bram[55637] = 243;
// bram[55638] = 231;
// bram[55639] = 215;
// bram[55640] = 196;
// bram[55641] = 175;
// bram[55642] = 151;
// bram[55643] = 127;
// bram[55644] = 102;
// bram[55645] = 79;
// bram[55646] = 57;
// bram[55647] = 38;
// bram[55648] = 22;
// bram[55649] = 10;
// bram[55650] = 2;
// bram[55651] = 0;
// bram[55652] = 1;
// bram[55653] = 8;
// bram[55654] = 19;
// bram[55655] = 34;
// bram[55656] = 52;
// bram[55657] = 73;
// bram[55658] = 97;
// bram[55659] = 121;
// bram[55660] = 145;
// bram[55661] = 169;
// bram[55662] = 191;
// bram[55663] = 211;
// bram[55664] = 228;
// bram[55665] = 241;
// bram[55666] = 249;
// bram[55667] = 253;
// bram[55668] = 252;
// bram[55669] = 247;
// bram[55670] = 237;
// bram[55671] = 223;
// bram[55672] = 205;
// bram[55673] = 185;
// bram[55674] = 162;
// bram[55675] = 138;
// bram[55676] = 113;
// bram[55677] = 89;
// bram[55678] = 66;
// bram[55679] = 46;
// bram[55680] = 29;
// bram[55681] = 15;
// bram[55682] = 5;
// bram[55683] = 0;
// bram[55684] = 0;
// bram[55685] = 4;
// bram[55686] = 13;
// bram[55687] = 26;
// bram[55688] = 43;
// bram[55689] = 63;
// bram[55690] = 86;
// bram[55691] = 110;
// bram[55692] = 134;
// bram[55693] = 159;
// bram[55694] = 182;
// bram[55695] = 203;
// bram[55696] = 221;
// bram[55697] = 235;
// bram[55698] = 246;
// bram[55699] = 252;
// bram[55700] = 253;
// bram[55701] = 250;
// bram[55702] = 242;
// bram[55703] = 230;
// bram[55704] = 214;
// bram[55705] = 194;
// bram[55706] = 172;
// bram[55707] = 149;
// bram[55708] = 124;
// bram[55709] = 100;
// bram[55710] = 77;
// bram[55711] = 55;
// bram[55712] = 36;
// bram[55713] = 21;
// bram[55714] = 9;
// bram[55715] = 2;
// bram[55716] = 0;
// bram[55717] = 2;
// bram[55718] = 9;
// bram[55719] = 20;
// bram[55720] = 35;
// bram[55721] = 54;
// bram[55722] = 75;
// bram[55723] = 99;
// bram[55724] = 123;
// bram[55725] = 148;
// bram[55726] = 171;
// bram[55727] = 193;
// bram[55728] = 213;
// bram[55729] = 229;
// bram[55730] = 242;
// bram[55731] = 250;
// bram[55732] = 253;
// bram[55733] = 252;
// bram[55734] = 246;
// bram[55735] = 236;
// bram[55736] = 221;
// bram[55737] = 204;
// bram[55738] = 183;
// bram[55739] = 160;
// bram[55740] = 135;
// bram[55741] = 111;
// bram[55742] = 87;
// bram[55743] = 64;
// bram[55744] = 44;
// bram[55745] = 27;
// bram[55746] = 14;
// bram[55747] = 5;
// bram[55748] = 0;
// bram[55749] = 0;
// bram[55750] = 5;
// bram[55751] = 14;
// bram[55752] = 28;
// bram[55753] = 45;
// bram[55754] = 65;
// bram[55755] = 88;
// bram[55756] = 112;
// bram[55757] = 137;
// bram[55758] = 161;
// bram[55759] = 184;
// bram[55760] = 204;
// bram[55761] = 222;
// bram[55762] = 236;
// bram[55763] = 247;
// bram[55764] = 252;
// bram[55765] = 253;
// bram[55766] = 250;
// bram[55767] = 241;
// bram[55768] = 229;
// bram[55769] = 212;
// bram[55770] = 192;
// bram[55771] = 170;
// bram[55772] = 147;
// bram[55773] = 122;
// bram[55774] = 98;
// bram[55775] = 74;
// bram[55776] = 53;
// bram[55777] = 35;
// bram[55778] = 19;
// bram[55779] = 8;
// bram[55780] = 2;
// bram[55781] = 0;
// bram[55782] = 2;
// bram[55783] = 10;
// bram[55784] = 21;
// bram[55785] = 37;
// bram[55786] = 56;
// bram[55787] = 77;
// bram[55788] = 101;
// bram[55789] = 125;
// bram[55790] = 150;
// bram[55791] = 173;
// bram[55792] = 195;
// bram[55793] = 214;
// bram[55794] = 230;
// bram[55795] = 243;
// bram[55796] = 250;
// bram[55797] = 253;
// bram[55798] = 252;
// bram[55799] = 246;
// bram[55800] = 235;
// bram[55801] = 220;
// bram[55802] = 202;
// bram[55803] = 181;
// bram[55804] = 158;
// bram[55805] = 133;
// bram[55806] = 109;
// bram[55807] = 85;
// bram[55808] = 63;
// bram[55809] = 43;
// bram[55810] = 26;
// bram[55811] = 13;
// bram[55812] = 4;
// bram[55813] = 0;
// bram[55814] = 0;
// bram[55815] = 6;
// bram[55816] = 15;
// bram[55817] = 29;
// bram[55818] = 47;
// bram[55819] = 67;
// bram[55820] = 90;
// bram[55821] = 114;
// bram[55822] = 139;
// bram[55823] = 163;
// bram[55824] = 186;
// bram[55825] = 206;
// bram[55826] = 224;
// bram[55827] = 238;
// bram[55828] = 247;
// bram[55829] = 253;
// bram[55830] = 253;
// bram[55831] = 249;
// bram[55832] = 240;
// bram[55833] = 227;
// bram[55834] = 210;
// bram[55835] = 191;
// bram[55836] = 168;
// bram[55837] = 144;
// bram[55838] = 120;
// bram[55839] = 96;
// bram[55840] = 72;
// bram[55841] = 51;
// bram[55842] = 33;
// bram[55843] = 18;
// bram[55844] = 7;
// bram[55845] = 1;
// bram[55846] = 0;
// bram[55847] = 3;
// bram[55848] = 10;
// bram[55849] = 23;
// bram[55850] = 38;
// bram[55851] = 58;
// bram[55852] = 80;
// bram[55853] = 103;
// bram[55854] = 128;
// bram[55855] = 152;
// bram[55856] = 175;
// bram[55857] = 197;
// bram[55858] = 216;
// bram[55859] = 232;
// bram[55860] = 243;
// bram[55861] = 251;
// bram[55862] = 253;
// bram[55863] = 251;
// bram[55864] = 245;
// bram[55865] = 234;
// bram[55866] = 218;
// bram[55867] = 200;
// bram[55868] = 179;
// bram[55869] = 155;
// bram[55870] = 131;
// bram[55871] = 106;
// bram[55872] = 83;
// bram[55873] = 61;
// bram[55874] = 41;
// bram[55875] = 24;
// bram[55876] = 12;
// bram[55877] = 3;
// bram[55878] = 0;
// bram[55879] = 1;
// bram[55880] = 6;
// bram[55881] = 17;
// bram[55882] = 31;
// bram[55883] = 49;
// bram[55884] = 69;
// bram[55885] = 92;
// bram[55886] = 116;
// bram[55887] = 141;
// bram[55888] = 165;
// bram[55889] = 188;
// bram[55890] = 208;
// bram[55891] = 225;
// bram[55892] = 239;
// bram[55893] = 248;
// bram[55894] = 253;
// bram[55895] = 253;
// bram[55896] = 248;
// bram[55897] = 239;
// bram[55898] = 226;
// bram[55899] = 209;
// bram[55900] = 189;
// bram[55901] = 166;
// bram[55902] = 142;
// bram[55903] = 118;
// bram[55904] = 93;
// bram[55905] = 70;
// bram[55906] = 50;
// bram[55907] = 32;
// bram[55908] = 17;
// bram[55909] = 7;
// bram[55910] = 1;
// bram[55911] = 0;
// bram[55912] = 3;
// bram[55913] = 11;
// bram[55914] = 24;
// bram[55915] = 40;
// bram[55916] = 60;
// bram[55917] = 82;
// bram[55918] = 105;
// bram[55919] = 130;
// bram[55920] = 154;
// bram[55921] = 178;
// bram[55922] = 199;
// bram[55923] = 218;
// bram[55924] = 233;
// bram[55925] = 244;
// bram[55926] = 251;
// bram[55927] = 253;
// bram[55928] = 251;
// bram[55929] = 244;
// bram[55930] = 232;
// bram[55931] = 217;
// bram[55932] = 198;
// bram[55933] = 177;
// bram[55934] = 153;
// bram[55935] = 129;
// bram[55936] = 104;
// bram[55937] = 81;
// bram[55938] = 59;
// bram[55939] = 39;
// bram[55940] = 23;
// bram[55941] = 11;
// bram[55942] = 3;
// bram[55943] = 0;
// bram[55944] = 1;
// bram[55945] = 7;
// bram[55946] = 18;
// bram[55947] = 32;
// bram[55948] = 50;
// bram[55949] = 71;
// bram[55950] = 94;
// bram[55951] = 119;
// bram[55952] = 143;
// bram[55953] = 167;
// bram[55954] = 190;
// bram[55955] = 210;
// bram[55956] = 226;
// bram[55957] = 240;
// bram[55958] = 249;
// bram[55959] = 253;
// bram[55960] = 253;
// bram[55961] = 248;
// bram[55962] = 238;
// bram[55963] = 224;
// bram[55964] = 207;
// bram[55965] = 187;
// bram[55966] = 164;
// bram[55967] = 140;
// bram[55968] = 115;
// bram[55969] = 91;
// bram[55970] = 68;
// bram[55971] = 48;
// bram[55972] = 30;
// bram[55973] = 16;
// bram[55974] = 6;
// bram[55975] = 1;
// bram[55976] = 0;
// bram[55977] = 4;
// bram[55978] = 12;
// bram[55979] = 25;
// bram[55980] = 42;
// bram[55981] = 62;
// bram[55982] = 84;
// bram[55983] = 108;
// bram[55984] = 132;
// bram[55985] = 156;
// bram[55986] = 180;
// bram[55987] = 201;
// bram[55988] = 219;
// bram[55989] = 234;
// bram[55990] = 245;
// bram[55991] = 252;
// bram[55992] = 253;
// bram[55993] = 251;
// bram[55994] = 243;
// bram[55995] = 231;
// bram[55996] = 215;
// bram[55997] = 196;
// bram[55998] = 174;
// bram[55999] = 151;
// bram[56000] = 127;
// bram[56001] = 152;
// bram[56002] = 177;
// bram[56003] = 200;
// bram[56004] = 219;
// bram[56005] = 235;
// bram[56006] = 246;
// bram[56007] = 252;
// bram[56008] = 253;
// bram[56009] = 249;
// bram[56010] = 239;
// bram[56011] = 225;
// bram[56012] = 206;
// bram[56013] = 184;
// bram[56014] = 160;
// bram[56015] = 134;
// bram[56016] = 108;
// bram[56017] = 83;
// bram[56018] = 60;
// bram[56019] = 39;
// bram[56020] = 22;
// bram[56021] = 9;
// bram[56022] = 2;
// bram[56023] = 0;
// bram[56024] = 2;
// bram[56025] = 11;
// bram[56026] = 24;
// bram[56027] = 41;
// bram[56028] = 62;
// bram[56029] = 86;
// bram[56030] = 111;
// bram[56031] = 137;
// bram[56032] = 163;
// bram[56033] = 187;
// bram[56034] = 208;
// bram[56035] = 226;
// bram[56036] = 240;
// bram[56037] = 249;
// bram[56038] = 253;
// bram[56039] = 252;
// bram[56040] = 245;
// bram[56041] = 234;
// bram[56042] = 217;
// bram[56043] = 198;
// bram[56044] = 175;
// bram[56045] = 150;
// bram[56046] = 124;
// bram[56047] = 98;
// bram[56048] = 73;
// bram[56049] = 51;
// bram[56050] = 32;
// bram[56051] = 16;
// bram[56052] = 6;
// bram[56053] = 0;
// bram[56054] = 0;
// bram[56055] = 5;
// bram[56056] = 15;
// bram[56057] = 30;
// bram[56058] = 49;
// bram[56059] = 71;
// bram[56060] = 96;
// bram[56061] = 122;
// bram[56062] = 148;
// bram[56063] = 173;
// bram[56064] = 196;
// bram[56065] = 216;
// bram[56066] = 233;
// bram[56067] = 245;
// bram[56068] = 252;
// bram[56069] = 253;
// bram[56070] = 250;
// bram[56071] = 241;
// bram[56072] = 228;
// bram[56073] = 210;
// bram[56074] = 188;
// bram[56075] = 165;
// bram[56076] = 139;
// bram[56077] = 113;
// bram[56078] = 88;
// bram[56079] = 64;
// bram[56080] = 43;
// bram[56081] = 25;
// bram[56082] = 11;
// bram[56083] = 3;
// bram[56084] = 0;
// bram[56085] = 2;
// bram[56086] = 9;
// bram[56087] = 21;
// bram[56088] = 38;
// bram[56089] = 58;
// bram[56090] = 81;
// bram[56091] = 106;
// bram[56092] = 132;
// bram[56093] = 158;
// bram[56094] = 182;
// bram[56095] = 205;
// bram[56096] = 223;
// bram[56097] = 238;
// bram[56098] = 248;
// bram[56099] = 253;
// bram[56100] = 253;
// bram[56101] = 247;
// bram[56102] = 236;
// bram[56103] = 221;
// bram[56104] = 201;
// bram[56105] = 179;
// bram[56106] = 154;
// bram[56107] = 128;
// bram[56108] = 103;
// bram[56109] = 78;
// bram[56110] = 55;
// bram[56111] = 35;
// bram[56112] = 19;
// bram[56113] = 7;
// bram[56114] = 1;
// bram[56115] = 0;
// bram[56116] = 4;
// bram[56117] = 13;
// bram[56118] = 27;
// bram[56119] = 45;
// bram[56120] = 67;
// bram[56121] = 91;
// bram[56122] = 117;
// bram[56123] = 143;
// bram[56124] = 168;
// bram[56125] = 192;
// bram[56126] = 213;
// bram[56127] = 230;
// bram[56128] = 243;
// bram[56129] = 251;
// bram[56130] = 253;
// bram[56131] = 251;
// bram[56132] = 243;
// bram[56133] = 230;
// bram[56134] = 213;
// bram[56135] = 193;
// bram[56136] = 169;
// bram[56137] = 144;
// bram[56138] = 118;
// bram[56139] = 92;
// bram[56140] = 68;
// bram[56141] = 46;
// bram[56142] = 28;
// bram[56143] = 14;
// bram[56144] = 4;
// bram[56145] = 0;
// bram[56146] = 1;
// bram[56147] = 7;
// bram[56148] = 18;
// bram[56149] = 34;
// bram[56150] = 54;
// bram[56151] = 77;
// bram[56152] = 102;
// bram[56153] = 127;
// bram[56154] = 153;
// bram[56155] = 178;
// bram[56156] = 201;
// bram[56157] = 220;
// bram[56158] = 236;
// bram[56159] = 247;
// bram[56160] = 252;
// bram[56161] = 253;
// bram[56162] = 248;
// bram[56163] = 239;
// bram[56164] = 224;
// bram[56165] = 205;
// bram[56166] = 183;
// bram[56167] = 159;
// bram[56168] = 133;
// bram[56169] = 107;
// bram[56170] = 82;
// bram[56171] = 59;
// bram[56172] = 38;
// bram[56173] = 21;
// bram[56174] = 9;
// bram[56175] = 2;
// bram[56176] = 0;
// bram[56177] = 3;
// bram[56178] = 11;
// bram[56179] = 24;
// bram[56180] = 42;
// bram[56181] = 63;
// bram[56182] = 87;
// bram[56183] = 112;
// bram[56184] = 138;
// bram[56185] = 164;
// bram[56186] = 188;
// bram[56187] = 209;
// bram[56188] = 227;
// bram[56189] = 241;
// bram[56190] = 250;
// bram[56191] = 253;
// bram[56192] = 252;
// bram[56193] = 245;
// bram[56194] = 233;
// bram[56195] = 217;
// bram[56196] = 197;
// bram[56197] = 174;
// bram[56198] = 149;
// bram[56199] = 123;
// bram[56200] = 97;
// bram[56201] = 72;
// bram[56202] = 50;
// bram[56203] = 31;
// bram[56204] = 16;
// bram[56205] = 5;
// bram[56206] = 0;
// bram[56207] = 0;
// bram[56208] = 5;
// bram[56209] = 16;
// bram[56210] = 31;
// bram[56211] = 50;
// bram[56212] = 72;
// bram[56213] = 97;
// bram[56214] = 123;
// bram[56215] = 149;
// bram[56216] = 174;
// bram[56217] = 197;
// bram[56218] = 217;
// bram[56219] = 233;
// bram[56220] = 245;
// bram[56221] = 252;
// bram[56222] = 253;
// bram[56223] = 250;
// bram[56224] = 241;
// bram[56225] = 227;
// bram[56226] = 209;
// bram[56227] = 188;
// bram[56228] = 164;
// bram[56229] = 138;
// bram[56230] = 112;
// bram[56231] = 87;
// bram[56232] = 63;
// bram[56233] = 42;
// bram[56234] = 24;
// bram[56235] = 11;
// bram[56236] = 3;
// bram[56237] = 0;
// bram[56238] = 2;
// bram[56239] = 9;
// bram[56240] = 21;
// bram[56241] = 38;
// bram[56242] = 59;
// bram[56243] = 82;
// bram[56244] = 107;
// bram[56245] = 133;
// bram[56246] = 159;
// bram[56247] = 183;
// bram[56248] = 205;
// bram[56249] = 224;
// bram[56250] = 239;
// bram[56251] = 248;
// bram[56252] = 253;
// bram[56253] = 253;
// bram[56254] = 247;
// bram[56255] = 236;
// bram[56256] = 220;
// bram[56257] = 201;
// bram[56258] = 178;
// bram[56259] = 153;
// bram[56260] = 127;
// bram[56261] = 102;
// bram[56262] = 77;
// bram[56263] = 54;
// bram[56264] = 34;
// bram[56265] = 18;
// bram[56266] = 7;
// bram[56267] = 1;
// bram[56268] = 0;
// bram[56269] = 4;
// bram[56270] = 14;
// bram[56271] = 28;
// bram[56272] = 46;
// bram[56273] = 68;
// bram[56274] = 92;
// bram[56275] = 118;
// bram[56276] = 144;
// bram[56277] = 169;
// bram[56278] = 193;
// bram[56279] = 213;
// bram[56280] = 230;
// bram[56281] = 243;
// bram[56282] = 251;
// bram[56283] = 253;
// bram[56284] = 251;
// bram[56285] = 243;
// bram[56286] = 230;
// bram[56287] = 213;
// bram[56288] = 192;
// bram[56289] = 168;
// bram[56290] = 143;
// bram[56291] = 117;
// bram[56292] = 91;
// bram[56293] = 67;
// bram[56294] = 45;
// bram[56295] = 27;
// bram[56296] = 13;
// bram[56297] = 4;
// bram[56298] = 0;
// bram[56299] = 1;
// bram[56300] = 7;
// bram[56301] = 19;
// bram[56302] = 35;
// bram[56303] = 55;
// bram[56304] = 78;
// bram[56305] = 102;
// bram[56306] = 128;
// bram[56307] = 154;
// bram[56308] = 179;
// bram[56309] = 201;
// bram[56310] = 221;
// bram[56311] = 236;
// bram[56312] = 247;
// bram[56313] = 253;
// bram[56314] = 253;
// bram[56315] = 248;
// bram[56316] = 238;
// bram[56317] = 223;
// bram[56318] = 205;
// bram[56319] = 183;
// bram[56320] = 158;
// bram[56321] = 132;
// bram[56322] = 106;
// bram[56323] = 81;
// bram[56324] = 58;
// bram[56325] = 38;
// bram[56326] = 21;
// bram[56327] = 9;
// bram[56328] = 2;
// bram[56329] = 0;
// bram[56330] = 3;
// bram[56331] = 11;
// bram[56332] = 25;
// bram[56333] = 42;
// bram[56334] = 64;
// bram[56335] = 87;
// bram[56336] = 113;
// bram[56337] = 139;
// bram[56338] = 165;
// bram[56339] = 188;
// bram[56340] = 210;
// bram[56341] = 228;
// bram[56342] = 241;
// bram[56343] = 250;
// bram[56344] = 253;
// bram[56345] = 252;
// bram[56346] = 245;
// bram[56347] = 233;
// bram[56348] = 216;
// bram[56349] = 196;
// bram[56350] = 173;
// bram[56351] = 148;
// bram[56352] = 122;
// bram[56353] = 96;
// bram[56354] = 71;
// bram[56355] = 49;
// bram[56356] = 30;
// bram[56357] = 15;
// bram[56358] = 5;
// bram[56359] = 0;
// bram[56360] = 0;
// bram[56361] = 6;
// bram[56362] = 16;
// bram[56363] = 32;
// bram[56364] = 51;
// bram[56365] = 73;
// bram[56366] = 98;
// bram[56367] = 124;
// bram[56368] = 150;
// bram[56369] = 175;
// bram[56370] = 197;
// bram[56371] = 217;
// bram[56372] = 234;
// bram[56373] = 245;
// bram[56374] = 252;
// bram[56375] = 253;
// bram[56376] = 249;
// bram[56377] = 240;
// bram[56378] = 226;
// bram[56379] = 208;
// bram[56380] = 187;
// bram[56381] = 163;
// bram[56382] = 137;
// bram[56383] = 111;
// bram[56384] = 86;
// bram[56385] = 62;
// bram[56386] = 41;
// bram[56387] = 24;
// bram[56388] = 11;
// bram[56389] = 2;
// bram[56390] = 0;
// bram[56391] = 2;
// bram[56392] = 9;
// bram[56393] = 22;
// bram[56394] = 39;
// bram[56395] = 60;
// bram[56396] = 83;
// bram[56397] = 108;
// bram[56398] = 134;
// bram[56399] = 160;
// bram[56400] = 184;
// bram[56401] = 206;
// bram[56402] = 225;
// bram[56403] = 239;
// bram[56404] = 249;
// bram[56405] = 253;
// bram[56406] = 252;
// bram[56407] = 246;
// bram[56408] = 235;
// bram[56409] = 220;
// bram[56410] = 200;
// bram[56411] = 177;
// bram[56412] = 152;
// bram[56413] = 127;
// bram[56414] = 101;
// bram[56415] = 76;
// bram[56416] = 53;
// bram[56417] = 34;
// bram[56418] = 18;
// bram[56419] = 7;
// bram[56420] = 1;
// bram[56421] = 0;
// bram[56422] = 4;
// bram[56423] = 14;
// bram[56424] = 28;
// bram[56425] = 47;
// bram[56426] = 69;
// bram[56427] = 93;
// bram[56428] = 119;
// bram[56429] = 145;
// bram[56430] = 170;
// bram[56431] = 193;
// bram[56432] = 214;
// bram[56433] = 231;
// bram[56434] = 243;
// bram[56435] = 251;
// bram[56436] = 253;
// bram[56437] = 251;
// bram[56438] = 242;
// bram[56439] = 229;
// bram[56440] = 212;
// bram[56441] = 191;
// bram[56442] = 167;
// bram[56443] = 142;
// bram[56444] = 116;
// bram[56445] = 90;
// bram[56446] = 66;
// bram[56447] = 45;
// bram[56448] = 27;
// bram[56449] = 13;
// bram[56450] = 4;
// bram[56451] = 0;
// bram[56452] = 1;
// bram[56453] = 8;
// bram[56454] = 19;
// bram[56455] = 35;
// bram[56456] = 55;
// bram[56457] = 78;
// bram[56458] = 103;
// bram[56459] = 129;
// bram[56460] = 155;
// bram[56461] = 180;
// bram[56462] = 202;
// bram[56463] = 221;
// bram[56464] = 237;
// bram[56465] = 247;
// bram[56466] = 253;
// bram[56467] = 253;
// bram[56468] = 248;
// bram[56469] = 238;
// bram[56470] = 223;
// bram[56471] = 204;
// bram[56472] = 182;
// bram[56473] = 157;
// bram[56474] = 131;
// bram[56475] = 105;
// bram[56476] = 80;
// bram[56477] = 57;
// bram[56478] = 37;
// bram[56479] = 20;
// bram[56480] = 8;
// bram[56481] = 1;
// bram[56482] = 0;
// bram[56483] = 3;
// bram[56484] = 12;
// bram[56485] = 25;
// bram[56486] = 43;
// bram[56487] = 64;
// bram[56488] = 88;
// bram[56489] = 114;
// bram[56490] = 140;
// bram[56491] = 165;
// bram[56492] = 189;
// bram[56493] = 210;
// bram[56494] = 228;
// bram[56495] = 242;
// bram[56496] = 250;
// bram[56497] = 253;
// bram[56498] = 251;
// bram[56499] = 244;
// bram[56500] = 232;
// bram[56501] = 215;
// bram[56502] = 195;
// bram[56503] = 172;
// bram[56504] = 147;
// bram[56505] = 121;
// bram[56506] = 95;
// bram[56507] = 71;
// bram[56508] = 49;
// bram[56509] = 30;
// bram[56510] = 15;
// bram[56511] = 5;
// bram[56512] = 0;
// bram[56513] = 0;
// bram[56514] = 6;
// bram[56515] = 17;
// bram[56516] = 32;
// bram[56517] = 51;
// bram[56518] = 74;
// bram[56519] = 99;
// bram[56520] = 125;
// bram[56521] = 150;
// bram[56522] = 175;
// bram[56523] = 198;
// bram[56524] = 218;
// bram[56525] = 234;
// bram[56526] = 246;
// bram[56527] = 252;
// bram[56528] = 253;
// bram[56529] = 249;
// bram[56530] = 240;
// bram[56531] = 226;
// bram[56532] = 208;
// bram[56533] = 186;
// bram[56534] = 162;
// bram[56535] = 136;
// bram[56536] = 110;
// bram[56537] = 85;
// bram[56538] = 61;
// bram[56539] = 40;
// bram[56540] = 23;
// bram[56541] = 10;
// bram[56542] = 2;
// bram[56543] = 0;
// bram[56544] = 2;
// bram[56545] = 10;
// bram[56546] = 23;
// bram[56547] = 40;
// bram[56548] = 60;
// bram[56549] = 84;
// bram[56550] = 109;
// bram[56551] = 135;
// bram[56552] = 161;
// bram[56553] = 185;
// bram[56554] = 207;
// bram[56555] = 225;
// bram[56556] = 239;
// bram[56557] = 249;
// bram[56558] = 253;
// bram[56559] = 252;
// bram[56560] = 246;
// bram[56561] = 235;
// bram[56562] = 219;
// bram[56563] = 199;
// bram[56564] = 176;
// bram[56565] = 152;
// bram[56566] = 126;
// bram[56567] = 100;
// bram[56568] = 75;
// bram[56569] = 52;
// bram[56570] = 33;
// bram[56571] = 17;
// bram[56572] = 6;
// bram[56573] = 1;
// bram[56574] = 0;
// bram[56575] = 5;
// bram[56576] = 14;
// bram[56577] = 29;
// bram[56578] = 48;
// bram[56579] = 70;
// bram[56580] = 94;
// bram[56581] = 120;
// bram[56582] = 146;
// bram[56583] = 171;
// bram[56584] = 194;
// bram[56585] = 215;
// bram[56586] = 231;
// bram[56587] = 244;
// bram[56588] = 251;
// bram[56589] = 253;
// bram[56590] = 250;
// bram[56591] = 242;
// bram[56592] = 229;
// bram[56593] = 211;
// bram[56594] = 190;
// bram[56595] = 166;
// bram[56596] = 141;
// bram[56597] = 115;
// bram[56598] = 89;
// bram[56599] = 65;
// bram[56600] = 44;
// bram[56601] = 26;
// bram[56602] = 12;
// bram[56603] = 3;
// bram[56604] = 0;
// bram[56605] = 1;
// bram[56606] = 8;
// bram[56607] = 20;
// bram[56608] = 36;
// bram[56609] = 56;
// bram[56610] = 79;
// bram[56611] = 104;
// bram[56612] = 130;
// bram[56613] = 156;
// bram[56614] = 181;
// bram[56615] = 203;
// bram[56616] = 222;
// bram[56617] = 237;
// bram[56618] = 247;
// bram[56619] = 253;
// bram[56620] = 253;
// bram[56621] = 248;
// bram[56622] = 237;
// bram[56623] = 222;
// bram[56624] = 203;
// bram[56625] = 181;
// bram[56626] = 156;
// bram[56627] = 130;
// bram[56628] = 104;
// bram[56629] = 79;
// bram[56630] = 56;
// bram[56631] = 36;
// bram[56632] = 20;
// bram[56633] = 8;
// bram[56634] = 1;
// bram[56635] = 0;
// bram[56636] = 3;
// bram[56637] = 12;
// bram[56638] = 26;
// bram[56639] = 44;
// bram[56640] = 65;
// bram[56641] = 89;
// bram[56642] = 115;
// bram[56643] = 141;
// bram[56644] = 166;
// bram[56645] = 190;
// bram[56646] = 211;
// bram[56647] = 229;
// bram[56648] = 242;
// bram[56649] = 250;
// bram[56650] = 253;
// bram[56651] = 251;
// bram[56652] = 244;
// bram[56653] = 232;
// bram[56654] = 215;
// bram[56655] = 194;
// bram[56656] = 171;
// bram[56657] = 146;
// bram[56658] = 120;
// bram[56659] = 94;
// bram[56660] = 70;
// bram[56661] = 48;
// bram[56662] = 29;
// bram[56663] = 15;
// bram[56664] = 5;
// bram[56665] = 0;
// bram[56666] = 0;
// bram[56667] = 6;
// bram[56668] = 17;
// bram[56669] = 33;
// bram[56670] = 52;
// bram[56671] = 75;
// bram[56672] = 100;
// bram[56673] = 125;
// bram[56674] = 151;
// bram[56675] = 176;
// bram[56676] = 199;
// bram[56677] = 219;
// bram[56678] = 235;
// bram[56679] = 246;
// bram[56680] = 252;
// bram[56681] = 253;
// bram[56682] = 249;
// bram[56683] = 239;
// bram[56684] = 225;
// bram[56685] = 207;
// bram[56686] = 185;
// bram[56687] = 161;
// bram[56688] = 135;
// bram[56689] = 109;
// bram[56690] = 84;
// bram[56691] = 60;
// bram[56692] = 40;
// bram[56693] = 23;
// bram[56694] = 10;
// bram[56695] = 2;
// bram[56696] = 0;
// bram[56697] = 2;
// bram[56698] = 10;
// bram[56699] = 23;
// bram[56700] = 40;
// bram[56701] = 61;
// bram[56702] = 85;
// bram[56703] = 110;
// bram[56704] = 136;
// bram[56705] = 162;
// bram[56706] = 186;
// bram[56707] = 207;
// bram[56708] = 226;
// bram[56709] = 240;
// bram[56710] = 249;
// bram[56711] = 253;
// bram[56712] = 252;
// bram[56713] = 246;
// bram[56714] = 234;
// bram[56715] = 218;
// bram[56716] = 198;
// bram[56717] = 176;
// bram[56718] = 151;
// bram[56719] = 125;
// bram[56720] = 99;
// bram[56721] = 74;
// bram[56722] = 52;
// bram[56723] = 32;
// bram[56724] = 17;
// bram[56725] = 6;
// bram[56726] = 0;
// bram[56727] = 0;
// bram[56728] = 5;
// bram[56729] = 15;
// bram[56730] = 30;
// bram[56731] = 48;
// bram[56732] = 70;
// bram[56733] = 95;
// bram[56734] = 121;
// bram[56735] = 147;
// bram[56736] = 172;
// bram[56737] = 195;
// bram[56738] = 215;
// bram[56739] = 232;
// bram[56740] = 244;
// bram[56741] = 251;
// bram[56742] = 253;
// bram[56743] = 250;
// bram[56744] = 242;
// bram[56745] = 228;
// bram[56746] = 211;
// bram[56747] = 189;
// bram[56748] = 166;
// bram[56749] = 140;
// bram[56750] = 114;
// bram[56751] = 89;
// bram[56752] = 65;
// bram[56753] = 43;
// bram[56754] = 25;
// bram[56755] = 12;
// bram[56756] = 3;
// bram[56757] = 0;
// bram[56758] = 1;
// bram[56759] = 8;
// bram[56760] = 20;
// bram[56761] = 37;
// bram[56762] = 57;
// bram[56763] = 80;
// bram[56764] = 105;
// bram[56765] = 131;
// bram[56766] = 157;
// bram[56767] = 182;
// bram[56768] = 204;
// bram[56769] = 223;
// bram[56770] = 238;
// bram[56771] = 248;
// bram[56772] = 253;
// bram[56773] = 253;
// bram[56774] = 247;
// bram[56775] = 237;
// bram[56776] = 221;
// bram[56777] = 202;
// bram[56778] = 180;
// bram[56779] = 155;
// bram[56780] = 129;
// bram[56781] = 104;
// bram[56782] = 79;
// bram[56783] = 56;
// bram[56784] = 36;
// bram[56785] = 19;
// bram[56786] = 8;
// bram[56787] = 1;
// bram[56788] = 0;
// bram[56789] = 4;
// bram[56790] = 13;
// bram[56791] = 27;
// bram[56792] = 45;
// bram[56793] = 66;
// bram[56794] = 90;
// bram[56795] = 116;
// bram[56796] = 142;
// bram[56797] = 167;
// bram[56798] = 191;
// bram[56799] = 212;
// bram[56800] = 229;
// bram[56801] = 242;
// bram[56802] = 251;
// bram[56803] = 253;
// bram[56804] = 251;
// bram[56805] = 244;
// bram[56806] = 231;
// bram[56807] = 214;
// bram[56808] = 194;
// bram[56809] = 170;
// bram[56810] = 145;
// bram[56811] = 119;
// bram[56812] = 93;
// bram[56813] = 69;
// bram[56814] = 47;
// bram[56815] = 28;
// bram[56816] = 14;
// bram[56817] = 4;
// bram[56818] = 0;
// bram[56819] = 1;
// bram[56820] = 7;
// bram[56821] = 18;
// bram[56822] = 33;
// bram[56823] = 53;
// bram[56824] = 76;
// bram[56825] = 101;
// bram[56826] = 126;
// bram[56827] = 152;
// bram[56828] = 177;
// bram[56829] = 200;
// bram[56830] = 219;
// bram[56831] = 235;
// bram[56832] = 246;
// bram[56833] = 252;
// bram[56834] = 253;
// bram[56835] = 249;
// bram[56836] = 239;
// bram[56837] = 225;
// bram[56838] = 206;
// bram[56839] = 184;
// bram[56840] = 160;
// bram[56841] = 134;
// bram[56842] = 108;
// bram[56843] = 83;
// bram[56844] = 60;
// bram[56845] = 39;
// bram[56846] = 22;
// bram[56847] = 10;
// bram[56848] = 2;
// bram[56849] = 0;
// bram[56850] = 2;
// bram[56851] = 11;
// bram[56852] = 24;
// bram[56853] = 41;
// bram[56854] = 62;
// bram[56855] = 86;
// bram[56856] = 111;
// bram[56857] = 137;
// bram[56858] = 163;
// bram[56859] = 187;
// bram[56860] = 208;
// bram[56861] = 226;
// bram[56862] = 240;
// bram[56863] = 249;
// bram[56864] = 253;
// bram[56865] = 252;
// bram[56866] = 245;
// bram[56867] = 234;
// bram[56868] = 218;
// bram[56869] = 198;
// bram[56870] = 175;
// bram[56871] = 150;
// bram[56872] = 124;
// bram[56873] = 98;
// bram[56874] = 73;
// bram[56875] = 51;
// bram[56876] = 32;
// bram[56877] = 16;
// bram[56878] = 6;
// bram[56879] = 0;
// bram[56880] = 0;
// bram[56881] = 5;
// bram[56882] = 15;
// bram[56883] = 30;
// bram[56884] = 49;
// bram[56885] = 71;
// bram[56886] = 96;
// bram[56887] = 122;
// bram[56888] = 148;
// bram[56889] = 173;
// bram[56890] = 196;
// bram[56891] = 216;
// bram[56892] = 233;
// bram[56893] = 245;
// bram[56894] = 252;
// bram[56895] = 253;
// bram[56896] = 250;
// bram[56897] = 241;
// bram[56898] = 228;
// bram[56899] = 210;
// bram[56900] = 189;
// bram[56901] = 165;
// bram[56902] = 139;
// bram[56903] = 113;
// bram[56904] = 88;
// bram[56905] = 64;
// bram[56906] = 43;
// bram[56907] = 25;
// bram[56908] = 12;
// bram[56909] = 3;
// bram[56910] = 0;
// bram[56911] = 2;
// bram[56912] = 9;
// bram[56913] = 21;
// bram[56914] = 37;
// bram[56915] = 58;
// bram[56916] = 81;
// bram[56917] = 106;
// bram[56918] = 132;
// bram[56919] = 158;
// bram[56920] = 182;
// bram[56921] = 204;
// bram[56922] = 223;
// bram[56923] = 238;
// bram[56924] = 248;
// bram[56925] = 253;
// bram[56926] = 253;
// bram[56927] = 247;
// bram[56928] = 236;
// bram[56929] = 221;
// bram[56930] = 202;
// bram[56931] = 179;
// bram[56932] = 154;
// bram[56933] = 129;
// bram[56934] = 103;
// bram[56935] = 78;
// bram[56936] = 55;
// bram[56937] = 35;
// bram[56938] = 19;
// bram[56939] = 7;
// bram[56940] = 1;
// bram[56941] = 0;
// bram[56942] = 4;
// bram[56943] = 13;
// bram[56944] = 27;
// bram[56945] = 45;
// bram[56946] = 67;
// bram[56947] = 91;
// bram[56948] = 117;
// bram[56949] = 143;
// bram[56950] = 168;
// bram[56951] = 192;
// bram[56952] = 213;
// bram[56953] = 230;
// bram[56954] = 243;
// bram[56955] = 251;
// bram[56956] = 253;
// bram[56957] = 251;
// bram[56958] = 243;
// bram[56959] = 230;
// bram[56960] = 213;
// bram[56961] = 193;
// bram[56962] = 169;
// bram[56963] = 144;
// bram[56964] = 118;
// bram[56965] = 92;
// bram[56966] = 68;
// bram[56967] = 46;
// bram[56968] = 28;
// bram[56969] = 14;
// bram[56970] = 4;
// bram[56971] = 0;
// bram[56972] = 1;
// bram[56973] = 7;
// bram[56974] = 18;
// bram[56975] = 34;
// bram[56976] = 54;
// bram[56977] = 77;
// bram[56978] = 101;
// bram[56979] = 127;
// bram[56980] = 153;
// bram[56981] = 178;
// bram[56982] = 201;
// bram[56983] = 220;
// bram[56984] = 236;
// bram[56985] = 247;
// bram[56986] = 252;
// bram[56987] = 253;
// bram[56988] = 248;
// bram[56989] = 239;
// bram[56990] = 224;
// bram[56991] = 205;
// bram[56992] = 183;
// bram[56993] = 159;
// bram[56994] = 133;
// bram[56995] = 107;
// bram[56996] = 82;
// bram[56997] = 59;
// bram[56998] = 38;
// bram[56999] = 22;
// bram[57000] = 9;
// bram[57001] = 2;
// bram[57002] = 0;
// bram[57003] = 3;
// bram[57004] = 11;
// bram[57005] = 24;
// bram[57006] = 42;
// bram[57007] = 63;
// bram[57008] = 86;
// bram[57009] = 112;
// bram[57010] = 138;
// bram[57011] = 164;
// bram[57012] = 188;
// bram[57013] = 209;
// bram[57014] = 227;
// bram[57015] = 241;
// bram[57016] = 250;
// bram[57017] = 253;
// bram[57018] = 252;
// bram[57019] = 245;
// bram[57020] = 233;
// bram[57021] = 217;
// bram[57022] = 197;
// bram[57023] = 174;
// bram[57024] = 149;
// bram[57025] = 123;
// bram[57026] = 97;
// bram[57027] = 72;
// bram[57028] = 50;
// bram[57029] = 31;
// bram[57030] = 16;
// bram[57031] = 6;
// bram[57032] = 0;
// bram[57033] = 0;
// bram[57034] = 5;
// bram[57035] = 16;
// bram[57036] = 31;
// bram[57037] = 50;
// bram[57038] = 72;
// bram[57039] = 97;
// bram[57040] = 123;
// bram[57041] = 148;
// bram[57042] = 174;
// bram[57043] = 197;
// bram[57044] = 217;
// bram[57045] = 233;
// bram[57046] = 245;
// bram[57047] = 252;
// bram[57048] = 253;
// bram[57049] = 250;
// bram[57050] = 241;
// bram[57051] = 227;
// bram[57052] = 209;
// bram[57053] = 188;
// bram[57054] = 164;
// bram[57055] = 138;
// bram[57056] = 112;
// bram[57057] = 87;
// bram[57058] = 63;
// bram[57059] = 42;
// bram[57060] = 24;
// bram[57061] = 11;
// bram[57062] = 3;
// bram[57063] = 0;
// bram[57064] = 2;
// bram[57065] = 9;
// bram[57066] = 21;
// bram[57067] = 38;
// bram[57068] = 59;
// bram[57069] = 82;
// bram[57070] = 107;
// bram[57071] = 133;
// bram[57072] = 159;
// bram[57073] = 183;
// bram[57074] = 205;
// bram[57075] = 224;
// bram[57076] = 238;
// bram[57077] = 248;
// bram[57078] = 253;
// bram[57079] = 253;
// bram[57080] = 247;
// bram[57081] = 236;
// bram[57082] = 220;
// bram[57083] = 201;
// bram[57084] = 178;
// bram[57085] = 153;
// bram[57086] = 128;
// bram[57087] = 102;
// bram[57088] = 77;
// bram[57089] = 54;
// bram[57090] = 34;
// bram[57091] = 18;
// bram[57092] = 7;
// bram[57093] = 1;
// bram[57094] = 0;
// bram[57095] = 4;
// bram[57096] = 14;
// bram[57097] = 28;
// bram[57098] = 46;
// bram[57099] = 68;
// bram[57100] = 92;
// bram[57101] = 118;
// bram[57102] = 144;
// bram[57103] = 169;
// bram[57104] = 193;
// bram[57105] = 213;
// bram[57106] = 230;
// bram[57107] = 243;
// bram[57108] = 251;
// bram[57109] = 253;
// bram[57110] = 251;
// bram[57111] = 243;
// bram[57112] = 230;
// bram[57113] = 213;
// bram[57114] = 192;
// bram[57115] = 168;
// bram[57116] = 143;
// bram[57117] = 117;
// bram[57118] = 91;
// bram[57119] = 67;
// bram[57120] = 46;
// bram[57121] = 27;
// bram[57122] = 13;
// bram[57123] = 4;
// bram[57124] = 0;
// bram[57125] = 1;
// bram[57126] = 7;
// bram[57127] = 19;
// bram[57128] = 35;
// bram[57129] = 55;
// bram[57130] = 77;
// bram[57131] = 102;
// bram[57132] = 128;
// bram[57133] = 154;
// bram[57134] = 179;
// bram[57135] = 201;
// bram[57136] = 221;
// bram[57137] = 236;
// bram[57138] = 247;
// bram[57139] = 253;
// bram[57140] = 253;
// bram[57141] = 248;
// bram[57142] = 238;
// bram[57143] = 223;
// bram[57144] = 205;
// bram[57145] = 183;
// bram[57146] = 158;
// bram[57147] = 132;
// bram[57148] = 106;
// bram[57149] = 81;
// bram[57150] = 58;
// bram[57151] = 38;
// bram[57152] = 21;
// bram[57153] = 9;
// bram[57154] = 2;
// bram[57155] = 0;
// bram[57156] = 3;
// bram[57157] = 11;
// bram[57158] = 25;
// bram[57159] = 42;
// bram[57160] = 64;
// bram[57161] = 87;
// bram[57162] = 113;
// bram[57163] = 139;
// bram[57164] = 164;
// bram[57165] = 188;
// bram[57166] = 210;
// bram[57167] = 227;
// bram[57168] = 241;
// bram[57169] = 250;
// bram[57170] = 253;
// bram[57171] = 252;
// bram[57172] = 245;
// bram[57173] = 233;
// bram[57174] = 216;
// bram[57175] = 196;
// bram[57176] = 173;
// bram[57177] = 148;
// bram[57178] = 122;
// bram[57179] = 96;
// bram[57180] = 72;
// bram[57181] = 49;
// bram[57182] = 30;
// bram[57183] = 15;
// bram[57184] = 5;
// bram[57185] = 0;
// bram[57186] = 0;
// bram[57187] = 6;
// bram[57188] = 16;
// bram[57189] = 31;
// bram[57190] = 51;
// bram[57191] = 73;
// bram[57192] = 98;
// bram[57193] = 123;
// bram[57194] = 149;
// bram[57195] = 174;
// bram[57196] = 197;
// bram[57197] = 217;
// bram[57198] = 234;
// bram[57199] = 245;
// bram[57200] = 252;
// bram[57201] = 253;
// bram[57202] = 249;
// bram[57203] = 240;
// bram[57204] = 226;
// bram[57205] = 208;
// bram[57206] = 187;
// bram[57207] = 163;
// bram[57208] = 137;
// bram[57209] = 111;
// bram[57210] = 86;
// bram[57211] = 62;
// bram[57212] = 41;
// bram[57213] = 24;
// bram[57214] = 11;
// bram[57215] = 3;
// bram[57216] = 0;
// bram[57217] = 2;
// bram[57218] = 9;
// bram[57219] = 22;
// bram[57220] = 39;
// bram[57221] = 59;
// bram[57222] = 83;
// bram[57223] = 108;
// bram[57224] = 134;
// bram[57225] = 160;
// bram[57226] = 184;
// bram[57227] = 206;
// bram[57228] = 224;
// bram[57229] = 239;
// bram[57230] = 249;
// bram[57231] = 253;
// bram[57232] = 252;
// bram[57233] = 246;
// bram[57234] = 235;
// bram[57235] = 220;
// bram[57236] = 200;
// bram[57237] = 177;
// bram[57238] = 153;
// bram[57239] = 127;
// bram[57240] = 101;
// bram[57241] = 76;
// bram[57242] = 53;
// bram[57243] = 34;
// bram[57244] = 18;
// bram[57245] = 7;
// bram[57246] = 1;
// bram[57247] = 0;
// bram[57248] = 4;
// bram[57249] = 14;
// bram[57250] = 28;
// bram[57251] = 47;
// bram[57252] = 69;
// bram[57253] = 93;
// bram[57254] = 119;
// bram[57255] = 145;
// bram[57256] = 170;
// bram[57257] = 193;
// bram[57258] = 214;
// bram[57259] = 231;
// bram[57260] = 243;
// bram[57261] = 251;
// bram[57262] = 253;
// bram[57263] = 251;
// bram[57264] = 242;
// bram[57265] = 229;
// bram[57266] = 212;
// bram[57267] = 191;
// bram[57268] = 167;
// bram[57269] = 142;
// bram[57270] = 116;
// bram[57271] = 90;
// bram[57272] = 66;
// bram[57273] = 45;
// bram[57274] = 27;
// bram[57275] = 13;
// bram[57276] = 4;
// bram[57277] = 0;
// bram[57278] = 1;
// bram[57279] = 8;
// bram[57280] = 19;
// bram[57281] = 35;
// bram[57282] = 55;
// bram[57283] = 78;
// bram[57284] = 103;
// bram[57285] = 129;
// bram[57286] = 155;
// bram[57287] = 180;
// bram[57288] = 202;
// bram[57289] = 221;
// bram[57290] = 237;
// bram[57291] = 247;
// bram[57292] = 253;
// bram[57293] = 253;
// bram[57294] = 248;
// bram[57295] = 238;
// bram[57296] = 223;
// bram[57297] = 204;
// bram[57298] = 182;
// bram[57299] = 157;
// bram[57300] = 131;
// bram[57301] = 106;
// bram[57302] = 80;
// bram[57303] = 57;
// bram[57304] = 37;
// bram[57305] = 20;
// bram[57306] = 8;
// bram[57307] = 1;
// bram[57308] = 0;
// bram[57309] = 3;
// bram[57310] = 12;
// bram[57311] = 25;
// bram[57312] = 43;
// bram[57313] = 64;
// bram[57314] = 88;
// bram[57315] = 114;
// bram[57316] = 140;
// bram[57317] = 165;
// bram[57318] = 189;
// bram[57319] = 210;
// bram[57320] = 228;
// bram[57321] = 241;
// bram[57322] = 250;
// bram[57323] = 253;
// bram[57324] = 252;
// bram[57325] = 244;
// bram[57326] = 232;
// bram[57327] = 216;
// bram[57328] = 195;
// bram[57329] = 172;
// bram[57330] = 147;
// bram[57331] = 121;
// bram[57332] = 95;
// bram[57333] = 71;
// bram[57334] = 49;
// bram[57335] = 30;
// bram[57336] = 15;
// bram[57337] = 5;
// bram[57338] = 0;
// bram[57339] = 0;
// bram[57340] = 6;
// bram[57341] = 17;
// bram[57342] = 32;
// bram[57343] = 51;
// bram[57344] = 74;
// bram[57345] = 99;
// bram[57346] = 124;
// bram[57347] = 150;
// bram[57348] = 175;
// bram[57349] = 198;
// bram[57350] = 218;
// bram[57351] = 234;
// bram[57352] = 246;
// bram[57353] = 252;
// bram[57354] = 253;
// bram[57355] = 249;
// bram[57356] = 240;
// bram[57357] = 226;
// bram[57358] = 208;
// bram[57359] = 186;
// bram[57360] = 162;
// bram[57361] = 136;
// bram[57362] = 110;
// bram[57363] = 85;
// bram[57364] = 61;
// bram[57365] = 40;
// bram[57366] = 23;
// bram[57367] = 10;
// bram[57368] = 2;
// bram[57369] = 0;
// bram[57370] = 2;
// bram[57371] = 10;
// bram[57372] = 22;
// bram[57373] = 40;
// bram[57374] = 60;
// bram[57375] = 84;
// bram[57376] = 109;
// bram[57377] = 135;
// bram[57378] = 161;
// bram[57379] = 185;
// bram[57380] = 207;
// bram[57381] = 225;
// bram[57382] = 239;
// bram[57383] = 249;
// bram[57384] = 253;
// bram[57385] = 252;
// bram[57386] = 246;
// bram[57387] = 235;
// bram[57388] = 219;
// bram[57389] = 199;
// bram[57390] = 176;
// bram[57391] = 152;
// bram[57392] = 126;
// bram[57393] = 100;
// bram[57394] = 75;
// bram[57395] = 52;
// bram[57396] = 33;
// bram[57397] = 17;
// bram[57398] = 6;
// bram[57399] = 1;
// bram[57400] = 0;
// bram[57401] = 5;
// bram[57402] = 14;
// bram[57403] = 29;
// bram[57404] = 48;
// bram[57405] = 70;
// bram[57406] = 94;
// bram[57407] = 120;
// bram[57408] = 146;
// bram[57409] = 171;
// bram[57410] = 194;
// bram[57411] = 215;
// bram[57412] = 231;
// bram[57413] = 244;
// bram[57414] = 251;
// bram[57415] = 253;
// bram[57416] = 250;
// bram[57417] = 242;
// bram[57418] = 229;
// bram[57419] = 211;
// bram[57420] = 190;
// bram[57421] = 167;
// bram[57422] = 141;
// bram[57423] = 115;
// bram[57424] = 90;
// bram[57425] = 66;
// bram[57426] = 44;
// bram[57427] = 26;
// bram[57428] = 12;
// bram[57429] = 3;
// bram[57430] = 0;
// bram[57431] = 1;
// bram[57432] = 8;
// bram[57433] = 20;
// bram[57434] = 36;
// bram[57435] = 56;
// bram[57436] = 79;
// bram[57437] = 104;
// bram[57438] = 130;
// bram[57439] = 156;
// bram[57440] = 181;
// bram[57441] = 203;
// bram[57442] = 222;
// bram[57443] = 237;
// bram[57444] = 247;
// bram[57445] = 253;
// bram[57446] = 253;
// bram[57447] = 248;
// bram[57448] = 237;
// bram[57449] = 222;
// bram[57450] = 203;
// bram[57451] = 181;
// bram[57452] = 156;
// bram[57453] = 131;
// bram[57454] = 105;
// bram[57455] = 80;
// bram[57456] = 56;
// bram[57457] = 36;
// bram[57458] = 20;
// bram[57459] = 8;
// bram[57460] = 1;
// bram[57461] = 0;
// bram[57462] = 3;
// bram[57463] = 12;
// bram[57464] = 26;
// bram[57465] = 44;
// bram[57466] = 65;
// bram[57467] = 89;
// bram[57468] = 115;
// bram[57469] = 141;
// bram[57470] = 166;
// bram[57471] = 190;
// bram[57472] = 211;
// bram[57473] = 229;
// bram[57474] = 242;
// bram[57475] = 250;
// bram[57476] = 253;
// bram[57477] = 251;
// bram[57478] = 244;
// bram[57479] = 232;
// bram[57480] = 215;
// bram[57481] = 194;
// bram[57482] = 171;
// bram[57483] = 146;
// bram[57484] = 120;
// bram[57485] = 94;
// bram[57486] = 70;
// bram[57487] = 48;
// bram[57488] = 29;
// bram[57489] = 15;
// bram[57490] = 5;
// bram[57491] = 0;
// bram[57492] = 0;
// bram[57493] = 6;
// bram[57494] = 17;
// bram[57495] = 33;
// bram[57496] = 52;
// bram[57497] = 75;
// bram[57498] = 99;
// bram[57499] = 125;
// bram[57500] = 151;
// bram[57501] = 176;
// bram[57502] = 199;
// bram[57503] = 219;
// bram[57504] = 235;
// bram[57505] = 246;
// bram[57506] = 252;
// bram[57507] = 253;
// bram[57508] = 249;
// bram[57509] = 239;
// bram[57510] = 225;
// bram[57511] = 207;
// bram[57512] = 185;
// bram[57513] = 161;
// bram[57514] = 135;
// bram[57515] = 109;
// bram[57516] = 84;
// bram[57517] = 61;
// bram[57518] = 40;
// bram[57519] = 23;
// bram[57520] = 10;
// bram[57521] = 2;
// bram[57522] = 0;
// bram[57523] = 2;
// bram[57524] = 10;
// bram[57525] = 23;
// bram[57526] = 40;
// bram[57527] = 61;
// bram[57528] = 85;
// bram[57529] = 110;
// bram[57530] = 136;
// bram[57531] = 162;
// bram[57532] = 186;
// bram[57533] = 207;
// bram[57534] = 226;
// bram[57535] = 240;
// bram[57536] = 249;
// bram[57537] = 253;
// bram[57538] = 252;
// bram[57539] = 246;
// bram[57540] = 234;
// bram[57541] = 218;
// bram[57542] = 198;
// bram[57543] = 176;
// bram[57544] = 151;
// bram[57545] = 125;
// bram[57546] = 99;
// bram[57547] = 74;
// bram[57548] = 52;
// bram[57549] = 32;
// bram[57550] = 17;
// bram[57551] = 6;
// bram[57552] = 0;
// bram[57553] = 0;
// bram[57554] = 5;
// bram[57555] = 15;
// bram[57556] = 30;
// bram[57557] = 48;
// bram[57558] = 70;
// bram[57559] = 95;
// bram[57560] = 121;
// bram[57561] = 147;
// bram[57562] = 172;
// bram[57563] = 195;
// bram[57564] = 215;
// bram[57565] = 232;
// bram[57566] = 244;
// bram[57567] = 251;
// bram[57568] = 253;
// bram[57569] = 250;
// bram[57570] = 242;
// bram[57571] = 228;
// bram[57572] = 211;
// bram[57573] = 189;
// bram[57574] = 166;
// bram[57575] = 140;
// bram[57576] = 114;
// bram[57577] = 89;
// bram[57578] = 65;
// bram[57579] = 43;
// bram[57580] = 26;
// bram[57581] = 12;
// bram[57582] = 3;
// bram[57583] = 0;
// bram[57584] = 1;
// bram[57585] = 8;
// bram[57586] = 20;
// bram[57587] = 37;
// bram[57588] = 57;
// bram[57589] = 80;
// bram[57590] = 105;
// bram[57591] = 131;
// bram[57592] = 157;
// bram[57593] = 181;
// bram[57594] = 204;
// bram[57595] = 223;
// bram[57596] = 238;
// bram[57597] = 248;
// bram[57598] = 253;
// bram[57599] = 253;
// bram[57600] = 247;
// bram[57601] = 237;
// bram[57602] = 222;
// bram[57603] = 202;
// bram[57604] = 180;
// bram[57605] = 155;
// bram[57606] = 130;
// bram[57607] = 104;
// bram[57608] = 79;
// bram[57609] = 56;
// bram[57610] = 36;
// bram[57611] = 19;
// bram[57612] = 8;
// bram[57613] = 1;
// bram[57614] = 0;
// bram[57615] = 4;
// bram[57616] = 13;
// bram[57617] = 26;
// bram[57618] = 45;
// bram[57619] = 66;
// bram[57620] = 90;
// bram[57621] = 116;
// bram[57622] = 142;
// bram[57623] = 167;
// bram[57624] = 191;
// bram[57625] = 212;
// bram[57626] = 229;
// bram[57627] = 242;
// bram[57628] = 250;
// bram[57629] = 253;
// bram[57630] = 251;
// bram[57631] = 244;
// bram[57632] = 231;
// bram[57633] = 214;
// bram[57634] = 194;
// bram[57635] = 170;
// bram[57636] = 145;
// bram[57637] = 119;
// bram[57638] = 93;
// bram[57639] = 69;
// bram[57640] = 47;
// bram[57641] = 29;
// bram[57642] = 14;
// bram[57643] = 4;
// bram[57644] = 0;
// bram[57645] = 1;
// bram[57646] = 7;
// bram[57647] = 18;
// bram[57648] = 33;
// bram[57649] = 53;
// bram[57650] = 76;
// bram[57651] = 100;
// bram[57652] = 126;
// bram[57653] = 152;
// bram[57654] = 177;
// bram[57655] = 200;
// bram[57656] = 219;
// bram[57657] = 235;
// bram[57658] = 246;
// bram[57659] = 252;
// bram[57660] = 253;
// bram[57661] = 249;
// bram[57662] = 239;
// bram[57663] = 225;
// bram[57664] = 206;
// bram[57665] = 184;
// bram[57666] = 160;
// bram[57667] = 134;
// bram[57668] = 108;
// bram[57669] = 83;
// bram[57670] = 60;
// bram[57671] = 39;
// bram[57672] = 22;
// bram[57673] = 10;
// bram[57674] = 2;
// bram[57675] = 0;
// bram[57676] = 2;
// bram[57677] = 11;
// bram[57678] = 24;
// bram[57679] = 41;
// bram[57680] = 62;
// bram[57681] = 86;
// bram[57682] = 111;
// bram[57683] = 137;
// bram[57684] = 163;
// bram[57685] = 187;
// bram[57686] = 208;
// bram[57687] = 226;
// bram[57688] = 240;
// bram[57689] = 249;
// bram[57690] = 253;
// bram[57691] = 252;
// bram[57692] = 245;
// bram[57693] = 234;
// bram[57694] = 218;
// bram[57695] = 198;
// bram[57696] = 175;
// bram[57697] = 150;
// bram[57698] = 124;
// bram[57699] = 98;
// bram[57700] = 73;
// bram[57701] = 51;
// bram[57702] = 32;
// bram[57703] = 16;
// bram[57704] = 6;
// bram[57705] = 0;
// bram[57706] = 0;
// bram[57707] = 5;
// bram[57708] = 15;
// bram[57709] = 30;
// bram[57710] = 49;
// bram[57711] = 71;
// bram[57712] = 96;
// bram[57713] = 121;
// bram[57714] = 147;
// bram[57715] = 173;
// bram[57716] = 196;
// bram[57717] = 216;
// bram[57718] = 232;
// bram[57719] = 245;
// bram[57720] = 252;
// bram[57721] = 253;
// bram[57722] = 250;
// bram[57723] = 241;
// bram[57724] = 228;
// bram[57725] = 210;
// bram[57726] = 189;
// bram[57727] = 165;
// bram[57728] = 139;
// bram[57729] = 113;
// bram[57730] = 88;
// bram[57731] = 64;
// bram[57732] = 43;
// bram[57733] = 25;
// bram[57734] = 12;
// bram[57735] = 3;
// bram[57736] = 0;
// bram[57737] = 1;
// bram[57738] = 9;
// bram[57739] = 21;
// bram[57740] = 37;
// bram[57741] = 58;
// bram[57742] = 81;
// bram[57743] = 106;
// bram[57744] = 132;
// bram[57745] = 158;
// bram[57746] = 182;
// bram[57747] = 204;
// bram[57748] = 223;
// bram[57749] = 238;
// bram[57750] = 248;
// bram[57751] = 253;
// bram[57752] = 253;
// bram[57753] = 247;
// bram[57754] = 236;
// bram[57755] = 221;
// bram[57756] = 202;
// bram[57757] = 179;
// bram[57758] = 154;
// bram[57759] = 129;
// bram[57760] = 103;
// bram[57761] = 78;
// bram[57762] = 55;
// bram[57763] = 35;
// bram[57764] = 19;
// bram[57765] = 7;
// bram[57766] = 1;
// bram[57767] = 0;
// bram[57768] = 4;
// bram[57769] = 13;
// bram[57770] = 27;
// bram[57771] = 45;
// bram[57772] = 67;
// bram[57773] = 91;
// bram[57774] = 117;
// bram[57775] = 143;
// bram[57776] = 168;
// bram[57777] = 192;
// bram[57778] = 212;
// bram[57779] = 230;
// bram[57780] = 243;
// bram[57781] = 251;
// bram[57782] = 253;
// bram[57783] = 251;
// bram[57784] = 243;
// bram[57785] = 231;
// bram[57786] = 214;
// bram[57787] = 193;
// bram[57788] = 169;
// bram[57789] = 144;
// bram[57790] = 118;
// bram[57791] = 92;
// bram[57792] = 68;
// bram[57793] = 46;
// bram[57794] = 28;
// bram[57795] = 14;
// bram[57796] = 4;
// bram[57797] = 0;
// bram[57798] = 1;
// bram[57799] = 7;
// bram[57800] = 18;
// bram[57801] = 34;
// bram[57802] = 54;
// bram[57803] = 76;
// bram[57804] = 101;
// bram[57805] = 127;
// bram[57806] = 153;
// bram[57807] = 178;
// bram[57808] = 201;
// bram[57809] = 220;
// bram[57810] = 236;
// bram[57811] = 247;
// bram[57812] = 252;
// bram[57813] = 253;
// bram[57814] = 248;
// bram[57815] = 239;
// bram[57816] = 224;
// bram[57817] = 205;
// bram[57818] = 184;
// bram[57819] = 159;
// bram[57820] = 133;
// bram[57821] = 107;
// bram[57822] = 82;
// bram[57823] = 59;
// bram[57824] = 38;
// bram[57825] = 22;
// bram[57826] = 9;
// bram[57827] = 2;
// bram[57828] = 0;
// bram[57829] = 3;
// bram[57830] = 11;
// bram[57831] = 24;
// bram[57832] = 42;
// bram[57833] = 63;
// bram[57834] = 86;
// bram[57835] = 112;
// bram[57836] = 138;
// bram[57837] = 163;
// bram[57838] = 187;
// bram[57839] = 209;
// bram[57840] = 227;
// bram[57841] = 241;
// bram[57842] = 250;
// bram[57843] = 253;
// bram[57844] = 252;
// bram[57845] = 245;
// bram[57846] = 233;
// bram[57847] = 217;
// bram[57848] = 197;
// bram[57849] = 174;
// bram[57850] = 149;
// bram[57851] = 123;
// bram[57852] = 97;
// bram[57853] = 72;
// bram[57854] = 50;
// bram[57855] = 31;
// bram[57856] = 16;
// bram[57857] = 6;
// bram[57858] = 0;
// bram[57859] = 0;
// bram[57860] = 5;
// bram[57861] = 16;
// bram[57862] = 31;
// bram[57863] = 50;
// bram[57864] = 72;
// bram[57865] = 97;
// bram[57866] = 122;
// bram[57867] = 148;
// bram[57868] = 173;
// bram[57869] = 197;
// bram[57870] = 217;
// bram[57871] = 233;
// bram[57872] = 245;
// bram[57873] = 252;
// bram[57874] = 253;
// bram[57875] = 250;
// bram[57876] = 241;
// bram[57877] = 227;
// bram[57878] = 209;
// bram[57879] = 188;
// bram[57880] = 164;
// bram[57881] = 138;
// bram[57882] = 112;
// bram[57883] = 87;
// bram[57884] = 63;
// bram[57885] = 42;
// bram[57886] = 24;
// bram[57887] = 11;
// bram[57888] = 3;
// bram[57889] = 0;
// bram[57890] = 2;
// bram[57891] = 9;
// bram[57892] = 21;
// bram[57893] = 38;
// bram[57894] = 59;
// bram[57895] = 82;
// bram[57896] = 107;
// bram[57897] = 133;
// bram[57898] = 159;
// bram[57899] = 183;
// bram[57900] = 205;
// bram[57901] = 224;
// bram[57902] = 238;
// bram[57903] = 248;
// bram[57904] = 253;
// bram[57905] = 253;
// bram[57906] = 247;
// bram[57907] = 236;
// bram[57908] = 220;
// bram[57909] = 201;
// bram[57910] = 178;
// bram[57911] = 154;
// bram[57912] = 128;
// bram[57913] = 102;
// bram[57914] = 77;
// bram[57915] = 54;
// bram[57916] = 34;
// bram[57917] = 18;
// bram[57918] = 7;
// bram[57919] = 1;
// bram[57920] = 0;
// bram[57921] = 4;
// bram[57922] = 13;
// bram[57923] = 28;
// bram[57924] = 46;
// bram[57925] = 68;
// bram[57926] = 92;
// bram[57927] = 118;
// bram[57928] = 144;
// bram[57929] = 169;
// bram[57930] = 192;
// bram[57931] = 213;
// bram[57932] = 230;
// bram[57933] = 243;
// bram[57934] = 251;
// bram[57935] = 253;
// bram[57936] = 251;
// bram[57937] = 243;
// bram[57938] = 230;
// bram[57939] = 213;
// bram[57940] = 192;
// bram[57941] = 168;
// bram[57942] = 143;
// bram[57943] = 117;
// bram[57944] = 91;
// bram[57945] = 67;
// bram[57946] = 46;
// bram[57947] = 27;
// bram[57948] = 13;
// bram[57949] = 4;
// bram[57950] = 0;
// bram[57951] = 1;
// bram[57952] = 7;
// bram[57953] = 19;
// bram[57954] = 35;
// bram[57955] = 54;
// bram[57956] = 77;
// bram[57957] = 102;
// bram[57958] = 128;
// bram[57959] = 154;
// bram[57960] = 179;
// bram[57961] = 201;
// bram[57962] = 221;
// bram[57963] = 236;
// bram[57964] = 247;
// bram[57965] = 253;
// bram[57966] = 253;
// bram[57967] = 248;
// bram[57968] = 238;
// bram[57969] = 223;
// bram[57970] = 205;
// bram[57971] = 183;
// bram[57972] = 158;
// bram[57973] = 133;
// bram[57974] = 107;
// bram[57975] = 81;
// bram[57976] = 58;
// bram[57977] = 38;
// bram[57978] = 21;
// bram[57979] = 9;
// bram[57980] = 2;
// bram[57981] = 0;
// bram[57982] = 3;
// bram[57983] = 11;
// bram[57984] = 25;
// bram[57985] = 42;
// bram[57986] = 63;
// bram[57987] = 87;
// bram[57988] = 113;
// bram[57989] = 139;
// bram[57990] = 164;
// bram[57991] = 188;
// bram[57992] = 210;
// bram[57993] = 227;
// bram[57994] = 241;
// bram[57995] = 250;
// bram[57996] = 253;
// bram[57997] = 252;
// bram[57998] = 245;
// bram[57999] = 233;
// bram[58000] = 216;
// bram[58001] = 196;
// bram[58002] = 173;
// bram[58003] = 148;
// bram[58004] = 122;
// bram[58005] = 96;
// bram[58006] = 72;
// bram[58007] = 49;
// bram[58008] = 30;
// bram[58009] = 16;
// bram[58010] = 5;
// bram[58011] = 0;
// bram[58012] = 0;
// bram[58013] = 6;
// bram[58014] = 16;
// bram[58015] = 31;
// bram[58016] = 51;
// bram[58017] = 73;
// bram[58018] = 98;
// bram[58019] = 123;
// bram[58020] = 149;
// bram[58021] = 174;
// bram[58022] = 197;
// bram[58023] = 217;
// bram[58024] = 234;
// bram[58025] = 245;
// bram[58026] = 252;
// bram[58027] = 253;
// bram[58028] = 249;
// bram[58029] = 240;
// bram[58030] = 227;
// bram[58031] = 208;
// bram[58032] = 187;
// bram[58033] = 163;
// bram[58034] = 137;
// bram[58035] = 111;
// bram[58036] = 86;
// bram[58037] = 62;
// bram[58038] = 41;
// bram[58039] = 24;
// bram[58040] = 11;
// bram[58041] = 3;
// bram[58042] = 0;
// bram[58043] = 2;
// bram[58044] = 9;
// bram[58045] = 22;
// bram[58046] = 39;
// bram[58047] = 59;
// bram[58048] = 83;
// bram[58049] = 108;
// bram[58050] = 134;
// bram[58051] = 160;
// bram[58052] = 184;
// bram[58053] = 206;
// bram[58054] = 224;
// bram[58055] = 239;
// bram[58056] = 249;
// bram[58057] = 253;
// bram[58058] = 252;
// bram[58059] = 246;
// bram[58060] = 235;
// bram[58061] = 220;
// bram[58062] = 200;
// bram[58063] = 177;
// bram[58064] = 153;
// bram[58065] = 127;
// bram[58066] = 101;
// bram[58067] = 76;
// bram[58068] = 53;
// bram[58069] = 34;
// bram[58070] = 18;
// bram[58071] = 7;
// bram[58072] = 1;
// bram[58073] = 0;
// bram[58074] = 4;
// bram[58075] = 14;
// bram[58076] = 28;
// bram[58077] = 47;
// bram[58078] = 69;
// bram[58079] = 93;
// bram[58080] = 119;
// bram[58081] = 145;
// bram[58082] = 170;
// bram[58083] = 193;
// bram[58084] = 214;
// bram[58085] = 231;
// bram[58086] = 243;
// bram[58087] = 251;
// bram[58088] = 253;
// bram[58089] = 251;
// bram[58090] = 242;
// bram[58091] = 229;
// bram[58092] = 212;
// bram[58093] = 191;
// bram[58094] = 168;
// bram[58095] = 142;
// bram[58096] = 116;
// bram[58097] = 91;
// bram[58098] = 66;
// bram[58099] = 45;
// bram[58100] = 27;
// bram[58101] = 13;
// bram[58102] = 4;
// bram[58103] = 0;
// bram[58104] = 1;
// bram[58105] = 8;
// bram[58106] = 19;
// bram[58107] = 35;
// bram[58108] = 55;
// bram[58109] = 78;
// bram[58110] = 103;
// bram[58111] = 129;
// bram[58112] = 155;
// bram[58113] = 180;
// bram[58114] = 202;
// bram[58115] = 221;
// bram[58116] = 237;
// bram[58117] = 247;
// bram[58118] = 253;
// bram[58119] = 253;
// bram[58120] = 248;
// bram[58121] = 238;
// bram[58122] = 223;
// bram[58123] = 204;
// bram[58124] = 182;
// bram[58125] = 157;
// bram[58126] = 132;
// bram[58127] = 106;
// bram[58128] = 80;
// bram[58129] = 57;
// bram[58130] = 37;
// bram[58131] = 21;
// bram[58132] = 8;
// bram[58133] = 1;
// bram[58134] = 0;
// bram[58135] = 3;
// bram[58136] = 12;
// bram[58137] = 25;
// bram[58138] = 43;
// bram[58139] = 64;
// bram[58140] = 88;
// bram[58141] = 114;
// bram[58142] = 140;
// bram[58143] = 165;
// bram[58144] = 189;
// bram[58145] = 210;
// bram[58146] = 228;
// bram[58147] = 241;
// bram[58148] = 250;
// bram[58149] = 253;
// bram[58150] = 252;
// bram[58151] = 244;
// bram[58152] = 232;
// bram[58153] = 216;
// bram[58154] = 195;
// bram[58155] = 172;
// bram[58156] = 147;
// bram[58157] = 121;
// bram[58158] = 95;
// bram[58159] = 71;
// bram[58160] = 49;
// bram[58161] = 30;
// bram[58162] = 15;
// bram[58163] = 5;
// bram[58164] = 0;
// bram[58165] = 0;
// bram[58166] = 6;
// bram[58167] = 17;
// bram[58168] = 32;
// bram[58169] = 51;
// bram[58170] = 74;
// bram[58171] = 98;
// bram[58172] = 124;
// bram[58173] = 150;
// bram[58174] = 175;
// bram[58175] = 198;
// bram[58176] = 218;
// bram[58177] = 234;
// bram[58178] = 246;
// bram[58179] = 252;
// bram[58180] = 253;
// bram[58181] = 249;
// bram[58182] = 240;
// bram[58183] = 226;
// bram[58184] = 208;
// bram[58185] = 186;
// bram[58186] = 162;
// bram[58187] = 136;
// bram[58188] = 110;
// bram[58189] = 85;
// bram[58190] = 61;
// bram[58191] = 41;
// bram[58192] = 23;
// bram[58193] = 10;
// bram[58194] = 2;
// bram[58195] = 0;
// bram[58196] = 2;
// bram[58197] = 10;
// bram[58198] = 22;
// bram[58199] = 39;
// bram[58200] = 60;
// bram[58201] = 84;
// bram[58202] = 109;
// bram[58203] = 135;
// bram[58204] = 161;
// bram[58205] = 185;
// bram[58206] = 207;
// bram[58207] = 225;
// bram[58208] = 239;
// bram[58209] = 249;
// bram[58210] = 253;
// bram[58211] = 252;
// bram[58212] = 246;
// bram[58213] = 235;
// bram[58214] = 219;
// bram[58215] = 199;
// bram[58216] = 177;
// bram[58217] = 152;
// bram[58218] = 126;
// bram[58219] = 100;
// bram[58220] = 75;
// bram[58221] = 53;
// bram[58222] = 33;
// bram[58223] = 17;
// bram[58224] = 6;
// bram[58225] = 1;
// bram[58226] = 0;
// bram[58227] = 5;
// bram[58228] = 14;
// bram[58229] = 29;
// bram[58230] = 47;
// bram[58231] = 69;
// bram[58232] = 94;
// bram[58233] = 119;
// bram[58234] = 145;
// bram[58235] = 171;
// bram[58236] = 194;
// bram[58237] = 215;
// bram[58238] = 231;
// bram[58239] = 244;
// bram[58240] = 251;
// bram[58241] = 253;
// bram[58242] = 250;
// bram[58243] = 242;
// bram[58244] = 229;
// bram[58245] = 211;
// bram[58246] = 190;
// bram[58247] = 167;
// bram[58248] = 141;
// bram[58249] = 115;
// bram[58250] = 90;
// bram[58251] = 66;
// bram[58252] = 44;
// bram[58253] = 26;
// bram[58254] = 12;
// bram[58255] = 3;
// bram[58256] = 0;
// bram[58257] = 1;
// bram[58258] = 8;
// bram[58259] = 20;
// bram[58260] = 36;
// bram[58261] = 56;
// bram[58262] = 79;
// bram[58263] = 104;
// bram[58264] = 130;
// bram[58265] = 156;
// bram[58266] = 180;
// bram[58267] = 203;
// bram[58268] = 222;
// bram[58269] = 237;
// bram[58270] = 247;
// bram[58271] = 253;
// bram[58272] = 253;
// bram[58273] = 248;
// bram[58274] = 237;
// bram[58275] = 222;
// bram[58276] = 203;
// bram[58277] = 181;
// bram[58278] = 156;
// bram[58279] = 131;
// bram[58280] = 105;
// bram[58281] = 80;
// bram[58282] = 57;
// bram[58283] = 36;
// bram[58284] = 20;
// bram[58285] = 8;
// bram[58286] = 1;
// bram[58287] = 0;
// bram[58288] = 3;
// bram[58289] = 12;
// bram[58290] = 26;
// bram[58291] = 44;
// bram[58292] = 65;
// bram[58293] = 89;
// bram[58294] = 115;
// bram[58295] = 141;
// bram[58296] = 166;
// bram[58297] = 190;
// bram[58298] = 211;
// bram[58299] = 229;
// bram[58300] = 242;
// bram[58301] = 250;
// bram[58302] = 253;
// bram[58303] = 251;
// bram[58304] = 244;
// bram[58305] = 232;
// bram[58306] = 215;
// bram[58307] = 195;
// bram[58308] = 171;
// bram[58309] = 146;
// bram[58310] = 120;
// bram[58311] = 94;
// bram[58312] = 70;
// bram[58313] = 48;
// bram[58314] = 29;
// bram[58315] = 15;
// bram[58316] = 5;
// bram[58317] = 0;
// bram[58318] = 0;
// bram[58319] = 6;
// bram[58320] = 17;
// bram[58321] = 33;
// bram[58322] = 52;
// bram[58323] = 75;
// bram[58324] = 99;
// bram[58325] = 125;
// bram[58326] = 151;
// bram[58327] = 176;
// bram[58328] = 199;
// bram[58329] = 219;
// bram[58330] = 235;
// bram[58331] = 246;
// bram[58332] = 252;
// bram[58333] = 253;
// bram[58334] = 249;
// bram[58335] = 240;
// bram[58336] = 225;
// bram[58337] = 207;
// bram[58338] = 185;
// bram[58339] = 161;
// bram[58340] = 135;
// bram[58341] = 109;
// bram[58342] = 84;
// bram[58343] = 61;
// bram[58344] = 40;
// bram[58345] = 23;
// bram[58346] = 10;
// bram[58347] = 2;
// bram[58348] = 0;
// bram[58349] = 2;
// bram[58350] = 10;
// bram[58351] = 23;
// bram[58352] = 40;
// bram[58353] = 61;
// bram[58354] = 85;
// bram[58355] = 110;
// bram[58356] = 136;
// bram[58357] = 162;
// bram[58358] = 186;
// bram[58359] = 207;
// bram[58360] = 226;
// bram[58361] = 240;
// bram[58362] = 249;
// bram[58363] = 253;
// bram[58364] = 252;
// bram[58365] = 246;
// bram[58366] = 234;
// bram[58367] = 218;
// bram[58368] = 199;
// bram[58369] = 176;
// bram[58370] = 151;
// bram[58371] = 125;
// bram[58372] = 99;
// bram[58373] = 74;
// bram[58374] = 52;
// bram[58375] = 32;
// bram[58376] = 17;
// bram[58377] = 6;
// bram[58378] = 0;
// bram[58379] = 0;
// bram[58380] = 5;
// bram[58381] = 15;
// bram[58382] = 29;
// bram[58383] = 48;
// bram[58384] = 70;
// bram[58385] = 95;
// bram[58386] = 120;
// bram[58387] = 146;
// bram[58388] = 172;
// bram[58389] = 195;
// bram[58390] = 215;
// bram[58391] = 232;
// bram[58392] = 244;
// bram[58393] = 251;
// bram[58394] = 253;
// bram[58395] = 250;
// bram[58396] = 242;
// bram[58397] = 228;
// bram[58398] = 211;
// bram[58399] = 190;
// bram[58400] = 166;
// bram[58401] = 140;
// bram[58402] = 114;
// bram[58403] = 89;
// bram[58404] = 65;
// bram[58405] = 43;
// bram[58406] = 26;
// bram[58407] = 12;
// bram[58408] = 3;
// bram[58409] = 0;
// bram[58410] = 1;
// bram[58411] = 8;
// bram[58412] = 20;
// bram[58413] = 37;
// bram[58414] = 57;
// bram[58415] = 80;
// bram[58416] = 105;
// bram[58417] = 131;
// bram[58418] = 157;
// bram[58419] = 181;
// bram[58420] = 204;
// bram[58421] = 223;
// bram[58422] = 237;
// bram[58423] = 248;
// bram[58424] = 253;
// bram[58425] = 253;
// bram[58426] = 247;
// bram[58427] = 237;
// bram[58428] = 222;
// bram[58429] = 202;
// bram[58430] = 180;
// bram[58431] = 156;
// bram[58432] = 130;
// bram[58433] = 104;
// bram[58434] = 79;
// bram[58435] = 56;
// bram[58436] = 36;
// bram[58437] = 20;
// bram[58438] = 8;
// bram[58439] = 1;
// bram[58440] = 0;
// bram[58441] = 4;
// bram[58442] = 13;
// bram[58443] = 26;
// bram[58444] = 44;
// bram[58445] = 66;
// bram[58446] = 90;
// bram[58447] = 116;
// bram[58448] = 142;
// bram[58449] = 167;
// bram[58450] = 191;
// bram[58451] = 212;
// bram[58452] = 229;
// bram[58453] = 242;
// bram[58454] = 250;
// bram[58455] = 253;
// bram[58456] = 251;
// bram[58457] = 244;
// bram[58458] = 231;
// bram[58459] = 214;
// bram[58460] = 194;
// bram[58461] = 170;
// bram[58462] = 145;
// bram[58463] = 119;
// bram[58464] = 93;
// bram[58465] = 69;
// bram[58466] = 47;
// bram[58467] = 29;
// bram[58468] = 14;
// bram[58469] = 4;
// bram[58470] = 0;
// bram[58471] = 1;
// bram[58472] = 7;
// bram[58473] = 18;
// bram[58474] = 33;
// bram[58475] = 53;
// bram[58476] = 76;
// bram[58477] = 100;
// bram[58478] = 126;
// bram[58479] = 152;
// bram[58480] = 177;
// bram[58481] = 200;
// bram[58482] = 219;
// bram[58483] = 235;
// bram[58484] = 246;
// bram[58485] = 252;
// bram[58486] = 253;
// bram[58487] = 249;
// bram[58488] = 239;
// bram[58489] = 225;
// bram[58490] = 206;
// bram[58491] = 184;
// bram[58492] = 160;
// bram[58493] = 135;
// bram[58494] = 109;
// bram[58495] = 83;
// bram[58496] = 60;
// bram[58497] = 39;
// bram[58498] = 22;
// bram[58499] = 10;
// bram[58500] = 2;
// bram[58501] = 0;
// bram[58502] = 2;
// bram[58503] = 11;
// bram[58504] = 24;
// bram[58505] = 41;
// bram[58506] = 62;
// bram[58507] = 85;
// bram[58508] = 111;
// bram[58509] = 137;
// bram[58510] = 162;
// bram[58511] = 186;
// bram[58512] = 208;
// bram[58513] = 226;
// bram[58514] = 240;
// bram[58515] = 249;
// bram[58516] = 253;
// bram[58517] = 252;
// bram[58518] = 245;
// bram[58519] = 234;
// bram[58520] = 218;
// bram[58521] = 198;
// bram[58522] = 175;
// bram[58523] = 150;
// bram[58524] = 124;
// bram[58525] = 98;
// bram[58526] = 73;
// bram[58527] = 51;
// bram[58528] = 32;
// bram[58529] = 17;
// bram[58530] = 6;
// bram[58531] = 0;
// bram[58532] = 0;
// bram[58533] = 5;
// bram[58534] = 15;
// bram[58535] = 30;
// bram[58536] = 49;
// bram[58537] = 71;
// bram[58538] = 96;
// bram[58539] = 121;
// bram[58540] = 147;
// bram[58541] = 172;
// bram[58542] = 196;
// bram[58543] = 216;
// bram[58544] = 232;
// bram[58545] = 244;
// bram[58546] = 252;
// bram[58547] = 253;
// bram[58548] = 250;
// bram[58549] = 241;
// bram[58550] = 228;
// bram[58551] = 210;
// bram[58552] = 189;
// bram[58553] = 165;
// bram[58554] = 139;
// bram[58555] = 113;
// bram[58556] = 88;
// bram[58557] = 64;
// bram[58558] = 43;
// bram[58559] = 25;
// bram[58560] = 12;
// bram[58561] = 3;
// bram[58562] = 0;
// bram[58563] = 1;
// bram[58564] = 9;
// bram[58565] = 21;
// bram[58566] = 37;
// bram[58567] = 58;
// bram[58568] = 81;
// bram[58569] = 106;
// bram[58570] = 132;
// bram[58571] = 158;
// bram[58572] = 182;
// bram[58573] = 204;
// bram[58574] = 223;
// bram[58575] = 238;
// bram[58576] = 248;
// bram[58577] = 253;
// bram[58578] = 253;
// bram[58579] = 247;
// bram[58580] = 236;
// bram[58581] = 221;
// bram[58582] = 202;
// bram[58583] = 179;
// bram[58584] = 155;
// bram[58585] = 129;
// bram[58586] = 103;
// bram[58587] = 78;
// bram[58588] = 55;
// bram[58589] = 35;
// bram[58590] = 19;
// bram[58591] = 7;
// bram[58592] = 1;
// bram[58593] = 0;
// bram[58594] = 4;
// bram[58595] = 13;
// bram[58596] = 27;
// bram[58597] = 45;
// bram[58598] = 67;
// bram[58599] = 91;
// bram[58600] = 117;
// bram[58601] = 143;
// bram[58602] = 168;
// bram[58603] = 192;
// bram[58604] = 212;
// bram[58605] = 230;
// bram[58606] = 243;
// bram[58607] = 251;
// bram[58608] = 253;
// bram[58609] = 251;
// bram[58610] = 243;
// bram[58611] = 231;
// bram[58612] = 214;
// bram[58613] = 193;
// bram[58614] = 169;
// bram[58615] = 144;
// bram[58616] = 118;
// bram[58617] = 92;
// bram[58618] = 68;
// bram[58619] = 46;
// bram[58620] = 28;
// bram[58621] = 14;
// bram[58622] = 4;
// bram[58623] = 0;
// bram[58624] = 1;
// bram[58625] = 7;
// bram[58626] = 18;
// bram[58627] = 34;
// bram[58628] = 54;
// bram[58629] = 76;
// bram[58630] = 101;
// bram[58631] = 127;
// bram[58632] = 153;
// bram[58633] = 178;
// bram[58634] = 200;
// bram[58635] = 220;
// bram[58636] = 236;
// bram[58637] = 247;
// bram[58638] = 252;
// bram[58639] = 253;
// bram[58640] = 248;
// bram[58641] = 239;
// bram[58642] = 224;
// bram[58643] = 206;
// bram[58644] = 184;
// bram[58645] = 159;
// bram[58646] = 134;
// bram[58647] = 108;
// bram[58648] = 82;
// bram[58649] = 59;
// bram[58650] = 38;
// bram[58651] = 22;
// bram[58652] = 9;
// bram[58653] = 2;
// bram[58654] = 0;
// bram[58655] = 3;
// bram[58656] = 11;
// bram[58657] = 24;
// bram[58658] = 42;
// bram[58659] = 63;
// bram[58660] = 86;
// bram[58661] = 112;
// bram[58662] = 138;
// bram[58663] = 163;
// bram[58664] = 187;
// bram[58665] = 209;
// bram[58666] = 227;
// bram[58667] = 241;
// bram[58668] = 250;
// bram[58669] = 253;
// bram[58670] = 252;
// bram[58671] = 245;
// bram[58672] = 233;
// bram[58673] = 217;
// bram[58674] = 197;
// bram[58675] = 174;
// bram[58676] = 149;
// bram[58677] = 123;
// bram[58678] = 97;
// bram[58679] = 73;
// bram[58680] = 50;
// bram[58681] = 31;
// bram[58682] = 16;
// bram[58683] = 6;
// bram[58684] = 0;
// bram[58685] = 0;
// bram[58686] = 5;
// bram[58687] = 16;
// bram[58688] = 31;
// bram[58689] = 50;
// bram[58690] = 72;
// bram[58691] = 97;
// bram[58692] = 122;
// bram[58693] = 148;
// bram[58694] = 173;
// bram[58695] = 196;
// bram[58696] = 217;
// bram[58697] = 233;
// bram[58698] = 245;
// bram[58699] = 252;
// bram[58700] = 253;
// bram[58701] = 250;
// bram[58702] = 241;
// bram[58703] = 227;
// bram[58704] = 209;
// bram[58705] = 188;
// bram[58706] = 164;
// bram[58707] = 138;
// bram[58708] = 112;
// bram[58709] = 87;
// bram[58710] = 63;
// bram[58711] = 42;
// bram[58712] = 24;
// bram[58713] = 11;
// bram[58714] = 3;
// bram[58715] = 0;
// bram[58716] = 2;
// bram[58717] = 9;
// bram[58718] = 21;
// bram[58719] = 38;
// bram[58720] = 58;
// bram[58721] = 82;
// bram[58722] = 107;
// bram[58723] = 133;
// bram[58724] = 159;
// bram[58725] = 183;
// bram[58726] = 205;
// bram[58727] = 224;
// bram[58728] = 238;
// bram[58729] = 248;
// bram[58730] = 253;
// bram[58731] = 253;
// bram[58732] = 247;
// bram[58733] = 236;
// bram[58734] = 220;
// bram[58735] = 201;
// bram[58736] = 178;
// bram[58737] = 154;
// bram[58738] = 128;
// bram[58739] = 102;
// bram[58740] = 77;
// bram[58741] = 54;
// bram[58742] = 34;
// bram[58743] = 19;
// bram[58744] = 7;
// bram[58745] = 1;
// bram[58746] = 0;
// bram[58747] = 4;
// bram[58748] = 13;
// bram[58749] = 28;
// bram[58750] = 46;
// bram[58751] = 68;
// bram[58752] = 92;
// bram[58753] = 117;
// bram[58754] = 144;
// bram[58755] = 169;
// bram[58756] = 192;
// bram[58757] = 213;
// bram[58758] = 230;
// bram[58759] = 243;
// bram[58760] = 251;
// bram[58761] = 253;
// bram[58762] = 251;
// bram[58763] = 243;
// bram[58764] = 230;
// bram[58765] = 213;
// bram[58766] = 192;
// bram[58767] = 169;
// bram[58768] = 143;
// bram[58769] = 117;
// bram[58770] = 92;
// bram[58771] = 67;
// bram[58772] = 46;
// bram[58773] = 27;
// bram[58774] = 13;
// bram[58775] = 4;
// bram[58776] = 0;
// bram[58777] = 1;
// bram[58778] = 7;
// bram[58779] = 19;
// bram[58780] = 35;
// bram[58781] = 54;
// bram[58782] = 77;
// bram[58783] = 102;
// bram[58784] = 128;
// bram[58785] = 154;
// bram[58786] = 179;
// bram[58787] = 201;
// bram[58788] = 221;
// bram[58789] = 236;
// bram[58790] = 247;
// bram[58791] = 253;
// bram[58792] = 253;
// bram[58793] = 248;
// bram[58794] = 238;
// bram[58795] = 224;
// bram[58796] = 205;
// bram[58797] = 183;
// bram[58798] = 158;
// bram[58799] = 133;
// bram[58800] = 107;
// bram[58801] = 81;
// bram[58802] = 58;
// bram[58803] = 38;
// bram[58804] = 21;
// bram[58805] = 9;
// bram[58806] = 2;
// bram[58807] = 0;
// bram[58808] = 3;
// bram[58809] = 11;
// bram[58810] = 25;
// bram[58811] = 42;
// bram[58812] = 63;
// bram[58813] = 87;
// bram[58814] = 113;
// bram[58815] = 139;
// bram[58816] = 164;
// bram[58817] = 188;
// bram[58818] = 210;
// bram[58819] = 227;
// bram[58820] = 241;
// bram[58821] = 250;
// bram[58822] = 253;
// bram[58823] = 252;
// bram[58824] = 245;
// bram[58825] = 233;
// bram[58826] = 216;
// bram[58827] = 196;
// bram[58828] = 173;
// bram[58829] = 148;
// bram[58830] = 122;
// bram[58831] = 96;
// bram[58832] = 72;
// bram[58833] = 49;
// bram[58834] = 31;
// bram[58835] = 16;
// bram[58836] = 5;
// bram[58837] = 0;
// bram[58838] = 0;
// bram[58839] = 6;
// bram[58840] = 16;
// bram[58841] = 31;
// bram[58842] = 50;
// bram[58843] = 73;
// bram[58844] = 97;
// bram[58845] = 123;
// bram[58846] = 149;
// bram[58847] = 174;
// bram[58848] = 197;
// bram[58849] = 217;
// bram[58850] = 233;
// bram[58851] = 245;
// bram[58852] = 252;
// bram[58853] = 253;
// bram[58854] = 249;
// bram[58855] = 240;
// bram[58856] = 227;
// bram[58857] = 209;
// bram[58858] = 187;
// bram[58859] = 163;
// bram[58860] = 137;
// bram[58861] = 111;
// bram[58862] = 86;
// bram[58863] = 62;
// bram[58864] = 41;
// bram[58865] = 24;
// bram[58866] = 11;
// bram[58867] = 3;
// bram[58868] = 0;
// bram[58869] = 2;
// bram[58870] = 9;
// bram[58871] = 22;
// bram[58872] = 39;
// bram[58873] = 59;
// bram[58874] = 83;
// bram[58875] = 108;
// bram[58876] = 134;
// bram[58877] = 160;
// bram[58878] = 184;
// bram[58879] = 206;
// bram[58880] = 224;
// bram[58881] = 239;
// bram[58882] = 249;
// bram[58883] = 253;
// bram[58884] = 252;
// bram[58885] = 246;
// bram[58886] = 235;
// bram[58887] = 220;
// bram[58888] = 200;
// bram[58889] = 178;
// bram[58890] = 153;
// bram[58891] = 127;
// bram[58892] = 101;
// bram[58893] = 76;
// bram[58894] = 53;
// bram[58895] = 34;
// bram[58896] = 18;
// bram[58897] = 7;
// bram[58898] = 1;
// bram[58899] = 0;
// bram[58900] = 4;
// bram[58901] = 14;
// bram[58902] = 28;
// bram[58903] = 47;
// bram[58904] = 68;
// bram[58905] = 93;
// bram[58906] = 118;
// bram[58907] = 144;
// bram[58908] = 170;
// bram[58909] = 193;
// bram[58910] = 214;
// bram[58911] = 231;
// bram[58912] = 243;
// bram[58913] = 251;
// bram[58914] = 253;
// bram[58915] = 251;
// bram[58916] = 242;
// bram[58917] = 230;
// bram[58918] = 212;
// bram[58919] = 191;
// bram[58920] = 168;
// bram[58921] = 142;
// bram[58922] = 116;
// bram[58923] = 91;
// bram[58924] = 67;
// bram[58925] = 45;
// bram[58926] = 27;
// bram[58927] = 13;
// bram[58928] = 4;
// bram[58929] = 0;
// bram[58930] = 1;
// bram[58931] = 8;
// bram[58932] = 19;
// bram[58933] = 35;
// bram[58934] = 55;
// bram[58935] = 78;
// bram[58936] = 103;
// bram[58937] = 129;
// bram[58938] = 155;
// bram[58939] = 180;
// bram[58940] = 202;
// bram[58941] = 221;
// bram[58942] = 236;
// bram[58943] = 247;
// bram[58944] = 253;
// bram[58945] = 253;
// bram[58946] = 248;
// bram[58947] = 238;
// bram[58948] = 223;
// bram[58949] = 204;
// bram[58950] = 182;
// bram[58951] = 157;
// bram[58952] = 132;
// bram[58953] = 106;
// bram[58954] = 81;
// bram[58955] = 57;
// bram[58956] = 37;
// bram[58957] = 21;
// bram[58958] = 9;
// bram[58959] = 1;
// bram[58960] = 0;
// bram[58961] = 3;
// bram[58962] = 12;
// bram[58963] = 25;
// bram[58964] = 43;
// bram[58965] = 64;
// bram[58966] = 88;
// bram[58967] = 114;
// bram[58968] = 140;
// bram[58969] = 165;
// bram[58970] = 189;
// bram[58971] = 210;
// bram[58972] = 228;
// bram[58973] = 241;
// bram[58974] = 250;
// bram[58975] = 253;
// bram[58976] = 252;
// bram[58977] = 244;
// bram[58978] = 232;
// bram[58979] = 216;
// bram[58980] = 195;
// bram[58981] = 172;
// bram[58982] = 147;
// bram[58983] = 121;
// bram[58984] = 95;
// bram[58985] = 71;
// bram[58986] = 49;
// bram[58987] = 30;
// bram[58988] = 15;
// bram[58989] = 5;
// bram[58990] = 0;
// bram[58991] = 0;
// bram[58992] = 6;
// bram[58993] = 17;
// bram[58994] = 32;
// bram[58995] = 51;
// bram[58996] = 74;
// bram[58997] = 98;
// bram[58998] = 124;
// bram[58999] = 150;
// bram[59000] = 175;
// bram[59001] = 198;
// bram[59002] = 218;
// bram[59003] = 234;
// bram[59004] = 246;
// bram[59005] = 252;
// bram[59006] = 253;
// bram[59007] = 249;
// bram[59008] = 240;
// bram[59009] = 226;
// bram[59010] = 208;
// bram[59011] = 186;
// bram[59012] = 162;
// bram[59013] = 137;
// bram[59014] = 110;
// bram[59015] = 85;
// bram[59016] = 62;
// bram[59017] = 41;
// bram[59018] = 23;
// bram[59019] = 10;
// bram[59020] = 2;
// bram[59021] = 0;
// bram[59022] = 2;
// bram[59023] = 10;
// bram[59024] = 22;
// bram[59025] = 39;
// bram[59026] = 60;
// bram[59027] = 84;
// bram[59028] = 109;
// bram[59029] = 135;
// bram[59030] = 160;
// bram[59031] = 185;
// bram[59032] = 207;
// bram[59033] = 225;
// bram[59034] = 239;
// bram[59035] = 249;
// bram[59036] = 253;
// bram[59037] = 252;
// bram[59038] = 246;
// bram[59039] = 235;
// bram[59040] = 219;
// bram[59041] = 199;
// bram[59042] = 177;
// bram[59043] = 152;
// bram[59044] = 126;
// bram[59045] = 100;
// bram[59046] = 75;
// bram[59047] = 53;
// bram[59048] = 33;
// bram[59049] = 18;
// bram[59050] = 7;
// bram[59051] = 1;
// bram[59052] = 0;
// bram[59053] = 5;
// bram[59054] = 14;
// bram[59055] = 29;
// bram[59056] = 47;
// bram[59057] = 69;
// bram[59058] = 94;
// bram[59059] = 119;
// bram[59060] = 145;
// bram[59061] = 171;
// bram[59062] = 194;
// bram[59063] = 214;
// bram[59064] = 231;
// bram[59065] = 244;
// bram[59066] = 251;
// bram[59067] = 253;
// bram[59068] = 250;
// bram[59069] = 242;
// bram[59070] = 229;
// bram[59071] = 211;
// bram[59072] = 190;
// bram[59073] = 167;
// bram[59074] = 141;
// bram[59075] = 115;
// bram[59076] = 90;
// bram[59077] = 66;
// bram[59078] = 44;
// bram[59079] = 26;
// bram[59080] = 12;
// bram[59081] = 3;
// bram[59082] = 0;
// bram[59083] = 1;
// bram[59084] = 8;
// bram[59085] = 20;
// bram[59086] = 36;
// bram[59087] = 56;
// bram[59088] = 79;
// bram[59089] = 104;
// bram[59090] = 130;
// bram[59091] = 156;
// bram[59092] = 180;
// bram[59093] = 203;
// bram[59094] = 222;
// bram[59095] = 237;
// bram[59096] = 247;
// bram[59097] = 253;
// bram[59098] = 253;
// bram[59099] = 248;
// bram[59100] = 237;
// bram[59101] = 222;
// bram[59102] = 203;
// bram[59103] = 181;
// bram[59104] = 157;
// bram[59105] = 131;
// bram[59106] = 105;
// bram[59107] = 80;
// bram[59108] = 57;
// bram[59109] = 36;
// bram[59110] = 20;
// bram[59111] = 8;
// bram[59112] = 1;
// bram[59113] = 0;
// bram[59114] = 3;
// bram[59115] = 12;
// bram[59116] = 26;
// bram[59117] = 44;
// bram[59118] = 65;
// bram[59119] = 89;
// bram[59120] = 115;
// bram[59121] = 141;
// bram[59122] = 166;
// bram[59123] = 190;
// bram[59124] = 211;
// bram[59125] = 229;
// bram[59126] = 242;
// bram[59127] = 250;
// bram[59128] = 253;
// bram[59129] = 251;
// bram[59130] = 244;
// bram[59131] = 232;
// bram[59132] = 215;
// bram[59133] = 195;
// bram[59134] = 171;
// bram[59135] = 146;
// bram[59136] = 120;
// bram[59137] = 94;
// bram[59138] = 70;
// bram[59139] = 48;
// bram[59140] = 29;
// bram[59141] = 15;
// bram[59142] = 5;
// bram[59143] = 0;
// bram[59144] = 0;
// bram[59145] = 6;
// bram[59146] = 17;
// bram[59147] = 33;
// bram[59148] = 52;
// bram[59149] = 75;
// bram[59150] = 99;
// bram[59151] = 125;
// bram[59152] = 151;
// bram[59153] = 176;
// bram[59154] = 199;
// bram[59155] = 219;
// bram[59156] = 234;
// bram[59157] = 246;
// bram[59158] = 252;
// bram[59159] = 253;
// bram[59160] = 249;
// bram[59161] = 240;
// bram[59162] = 225;
// bram[59163] = 207;
// bram[59164] = 185;
// bram[59165] = 161;
// bram[59166] = 136;
// bram[59167] = 110;
// bram[59168] = 84;
// bram[59169] = 61;
// bram[59170] = 40;
// bram[59171] = 23;
// bram[59172] = 10;
// bram[59173] = 2;
// bram[59174] = 0;
// bram[59175] = 2;
// bram[59176] = 10;
// bram[59177] = 23;
// bram[59178] = 40;
// bram[59179] = 61;
// bram[59180] = 84;
// bram[59181] = 110;
// bram[59182] = 136;
// bram[59183] = 161;
// bram[59184] = 186;
// bram[59185] = 207;
// bram[59186] = 226;
// bram[59187] = 240;
// bram[59188] = 249;
// bram[59189] = 253;
// bram[59190] = 252;
// bram[59191] = 246;
// bram[59192] = 234;
// bram[59193] = 218;
// bram[59194] = 199;
// bram[59195] = 176;
// bram[59196] = 151;
// bram[59197] = 125;
// bram[59198] = 99;
// bram[59199] = 74;
// bram[59200] = 52;
// bram[59201] = 32;
// bram[59202] = 17;
// bram[59203] = 6;
// bram[59204] = 0;
// bram[59205] = 0;
// bram[59206] = 5;
// bram[59207] = 15;
// bram[59208] = 29;
// bram[59209] = 48;
// bram[59210] = 70;
// bram[59211] = 95;
// bram[59212] = 120;
// bram[59213] = 146;
// bram[59214] = 171;
// bram[59215] = 195;
// bram[59216] = 215;
// bram[59217] = 232;
// bram[59218] = 244;
// bram[59219] = 251;
// bram[59220] = 253;
// bram[59221] = 250;
// bram[59222] = 242;
// bram[59223] = 228;
// bram[59224] = 211;
// bram[59225] = 190;
// bram[59226] = 166;
// bram[59227] = 140;
// bram[59228] = 114;
// bram[59229] = 89;
// bram[59230] = 65;
// bram[59231] = 44;
// bram[59232] = 26;
// bram[59233] = 12;
// bram[59234] = 3;
// bram[59235] = 0;
// bram[59236] = 1;
// bram[59237] = 8;
// bram[59238] = 20;
// bram[59239] = 37;
// bram[59240] = 57;
// bram[59241] = 80;
// bram[59242] = 105;
// bram[59243] = 131;
// bram[59244] = 157;
// bram[59245] = 181;
// bram[59246] = 203;
// bram[59247] = 222;
// bram[59248] = 237;
// bram[59249] = 248;
// bram[59250] = 253;
// bram[59251] = 253;
// bram[59252] = 247;
// bram[59253] = 237;
// bram[59254] = 222;
// bram[59255] = 203;
// bram[59256] = 180;
// bram[59257] = 156;
// bram[59258] = 130;
// bram[59259] = 104;
// bram[59260] = 79;
// bram[59261] = 56;
// bram[59262] = 36;
// bram[59263] = 20;
// bram[59264] = 8;
// bram[59265] = 1;
// bram[59266] = 0;
// bram[59267] = 4;
// bram[59268] = 13;
// bram[59269] = 26;
// bram[59270] = 44;
// bram[59271] = 66;
// bram[59272] = 90;
// bram[59273] = 115;
// bram[59274] = 142;
// bram[59275] = 167;
// bram[59276] = 191;
// bram[59277] = 212;
// bram[59278] = 229;
// bram[59279] = 242;
// bram[59280] = 250;
// bram[59281] = 253;
// bram[59282] = 251;
// bram[59283] = 244;
// bram[59284] = 231;
// bram[59285] = 214;
// bram[59286] = 194;
// bram[59287] = 170;
// bram[59288] = 145;
// bram[59289] = 119;
// bram[59290] = 93;
// bram[59291] = 69;
// bram[59292] = 47;
// bram[59293] = 29;
// bram[59294] = 14;
// bram[59295] = 4;
// bram[59296] = 0;
// bram[59297] = 1;
// bram[59298] = 7;
// bram[59299] = 18;
// bram[59300] = 33;
// bram[59301] = 53;
// bram[59302] = 75;
// bram[59303] = 100;
// bram[59304] = 126;
// bram[59305] = 152;
// bram[59306] = 177;
// bram[59307] = 200;
// bram[59308] = 219;
// bram[59309] = 235;
// bram[59310] = 246;
// bram[59311] = 252;
// bram[59312] = 253;
// bram[59313] = 249;
// bram[59314] = 239;
// bram[59315] = 225;
// bram[59316] = 206;
// bram[59317] = 185;
// bram[59318] = 160;
// bram[59319] = 135;
// bram[59320] = 109;
// bram[59321] = 83;
// bram[59322] = 60;
// bram[59323] = 39;
// bram[59324] = 22;
// bram[59325] = 10;
// bram[59326] = 2;
// bram[59327] = 0;
// bram[59328] = 2;
// bram[59329] = 10;
// bram[59330] = 23;
// bram[59331] = 41;
// bram[59332] = 62;
// bram[59333] = 85;
// bram[59334] = 111;
// bram[59335] = 137;
// bram[59336] = 162;
// bram[59337] = 186;
// bram[59338] = 208;
// bram[59339] = 226;
// bram[59340] = 240;
// bram[59341] = 249;
// bram[59342] = 253;
// bram[59343] = 252;
// bram[59344] = 245;
// bram[59345] = 234;
// bram[59346] = 218;
// bram[59347] = 198;
// bram[59348] = 175;
// bram[59349] = 150;
// bram[59350] = 124;
// bram[59351] = 98;
// bram[59352] = 74;
// bram[59353] = 51;
// bram[59354] = 32;
// bram[59355] = 17;
// bram[59356] = 6;
// bram[59357] = 0;
// bram[59358] = 0;
// bram[59359] = 5;
// bram[59360] = 15;
// bram[59361] = 30;
// bram[59362] = 49;
// bram[59363] = 71;
// bram[59364] = 95;
// bram[59365] = 121;
// bram[59366] = 147;
// bram[59367] = 172;
// bram[59368] = 196;
// bram[59369] = 216;
// bram[59370] = 232;
// bram[59371] = 244;
// bram[59372] = 252;
// bram[59373] = 253;
// bram[59374] = 250;
// bram[59375] = 241;
// bram[59376] = 228;
// bram[59377] = 210;
// bram[59378] = 189;
// bram[59379] = 165;
// bram[59380] = 139;
// bram[59381] = 113;
// bram[59382] = 88;
// bram[59383] = 64;
// bram[59384] = 43;
// bram[59385] = 25;
// bram[59386] = 12;
// bram[59387] = 3;
// bram[59388] = 0;
// bram[59389] = 1;
// bram[59390] = 9;
// bram[59391] = 21;
// bram[59392] = 37;
// bram[59393] = 58;
// bram[59394] = 81;
// bram[59395] = 106;
// bram[59396] = 132;
// bram[59397] = 158;
// bram[59398] = 182;
// bram[59399] = 204;
// bram[59400] = 223;
// bram[59401] = 238;
// bram[59402] = 248;
// bram[59403] = 253;
// bram[59404] = 253;
// bram[59405] = 247;
// bram[59406] = 236;
// bram[59407] = 221;
// bram[59408] = 202;
// bram[59409] = 179;
// bram[59410] = 155;
// bram[59411] = 129;
// bram[59412] = 103;
// bram[59413] = 78;
// bram[59414] = 55;
// bram[59415] = 35;
// bram[59416] = 19;
// bram[59417] = 8;
// bram[59418] = 1;
// bram[59419] = 0;
// bram[59420] = 4;
// bram[59421] = 13;
// bram[59422] = 27;
// bram[59423] = 45;
// bram[59424] = 67;
// bram[59425] = 91;
// bram[59426] = 116;
// bram[59427] = 142;
// bram[59428] = 168;
// bram[59429] = 191;
// bram[59430] = 212;
// bram[59431] = 230;
// bram[59432] = 243;
// bram[59433] = 251;
// bram[59434] = 253;
// bram[59435] = 251;
// bram[59436] = 243;
// bram[59437] = 231;
// bram[59438] = 214;
// bram[59439] = 193;
// bram[59440] = 170;
// bram[59441] = 144;
// bram[59442] = 118;
// bram[59443] = 93;
// bram[59444] = 68;
// bram[59445] = 47;
// bram[59446] = 28;
// bram[59447] = 14;
// bram[59448] = 4;
// bram[59449] = 0;
// bram[59450] = 1;
// bram[59451] = 7;
// bram[59452] = 18;
// bram[59453] = 34;
// bram[59454] = 54;
// bram[59455] = 76;
// bram[59456] = 101;
// bram[59457] = 127;
// bram[59458] = 153;
// bram[59459] = 178;
// bram[59460] = 200;
// bram[59461] = 220;
// bram[59462] = 235;
// bram[59463] = 246;
// bram[59464] = 252;
// bram[59465] = 253;
// bram[59466] = 248;
// bram[59467] = 239;
// bram[59468] = 224;
// bram[59469] = 206;
// bram[59470] = 184;
// bram[59471] = 159;
// bram[59472] = 134;
// bram[59473] = 108;
// bram[59474] = 82;
// bram[59475] = 59;
// bram[59476] = 39;
// bram[59477] = 22;
// bram[59478] = 9;
// bram[59479] = 2;
// bram[59480] = 0;
// bram[59481] = 3;
// bram[59482] = 11;
// bram[59483] = 24;
// bram[59484] = 41;
// bram[59485] = 62;
// bram[59486] = 86;
// bram[59487] = 112;
// bram[59488] = 138;
// bram[59489] = 163;
// bram[59490] = 187;
// bram[59491] = 209;
// bram[59492] = 227;
// bram[59493] = 241;
// bram[59494] = 250;
// bram[59495] = 253;
// bram[59496] = 252;
// bram[59497] = 245;
// bram[59498] = 233;
// bram[59499] = 217;
// bram[59500] = 197;
// bram[59501] = 174;
// bram[59502] = 149;
// bram[59503] = 123;
// bram[59504] = 97;
// bram[59505] = 73;
// bram[59506] = 50;
// bram[59507] = 31;
// bram[59508] = 16;
// bram[59509] = 6;
// bram[59510] = 0;
// bram[59511] = 0;
// bram[59512] = 5;
// bram[59513] = 16;
// bram[59514] = 31;
// bram[59515] = 50;
// bram[59516] = 72;
// bram[59517] = 96;
// bram[59518] = 122;
// bram[59519] = 148;
// bram[59520] = 173;
// bram[59521] = 196;
// bram[59522] = 217;
// bram[59523] = 233;
// bram[59524] = 245;
// bram[59525] = 252;
// bram[59526] = 253;
// bram[59527] = 250;
// bram[59528] = 241;
// bram[59529] = 227;
// bram[59530] = 209;
// bram[59531] = 188;
// bram[59532] = 164;
// bram[59533] = 139;
// bram[59534] = 112;
// bram[59535] = 87;
// bram[59536] = 63;
// bram[59537] = 42;
// bram[59538] = 25;
// bram[59539] = 11;
// bram[59540] = 3;
// bram[59541] = 0;
// bram[59542] = 2;
// bram[59543] = 9;
// bram[59544] = 21;
// bram[59545] = 38;
// bram[59546] = 58;
// bram[59547] = 82;
// bram[59548] = 107;
// bram[59549] = 133;
// bram[59550] = 159;
// bram[59551] = 183;
// bram[59552] = 205;
// bram[59553] = 224;
// bram[59554] = 238;
// bram[59555] = 248;
// bram[59556] = 253;
// bram[59557] = 253;
// bram[59558] = 247;
// bram[59559] = 236;
// bram[59560] = 220;
// bram[59561] = 201;
// bram[59562] = 178;
// bram[59563] = 154;
// bram[59564] = 128;
// bram[59565] = 102;
// bram[59566] = 77;
// bram[59567] = 54;
// bram[59568] = 34;
// bram[59569] = 19;
// bram[59570] = 7;
// bram[59571] = 1;
// bram[59572] = 0;
// bram[59573] = 4;
// bram[59574] = 13;
// bram[59575] = 28;
// bram[59576] = 46;
// bram[59577] = 68;
// bram[59578] = 92;
// bram[59579] = 117;
// bram[59580] = 143;
// bram[59581] = 169;
// bram[59582] = 192;
// bram[59583] = 213;
// bram[59584] = 230;
// bram[59585] = 243;
// bram[59586] = 251;
// bram[59587] = 253;
// bram[59588] = 251;
// bram[59589] = 243;
// bram[59590] = 230;
// bram[59591] = 213;
// bram[59592] = 192;
// bram[59593] = 169;
// bram[59594] = 143;
// bram[59595] = 117;
// bram[59596] = 92;
// bram[59597] = 67;
// bram[59598] = 46;
// bram[59599] = 27;
// bram[59600] = 13;
// bram[59601] = 4;
// bram[59602] = 0;
// bram[59603] = 1;
// bram[59604] = 7;
// bram[59605] = 19;
// bram[59606] = 35;
// bram[59607] = 54;
// bram[59608] = 77;
// bram[59609] = 102;
// bram[59610] = 128;
// bram[59611] = 154;
// bram[59612] = 179;
// bram[59613] = 201;
// bram[59614] = 221;
// bram[59615] = 236;
// bram[59616] = 247;
// bram[59617] = 253;
// bram[59618] = 253;
// bram[59619] = 248;
// bram[59620] = 238;
// bram[59621] = 224;
// bram[59622] = 205;
// bram[59623] = 183;
// bram[59624] = 158;
// bram[59625] = 133;
// bram[59626] = 107;
// bram[59627] = 82;
// bram[59628] = 58;
// bram[59629] = 38;
// bram[59630] = 21;
// bram[59631] = 9;
// bram[59632] = 2;
// bram[59633] = 0;
// bram[59634] = 3;
// bram[59635] = 11;
// bram[59636] = 25;
// bram[59637] = 42;
// bram[59638] = 63;
// bram[59639] = 87;
// bram[59640] = 113;
// bram[59641] = 139;
// bram[59642] = 164;
// bram[59643] = 188;
// bram[59644] = 209;
// bram[59645] = 227;
// bram[59646] = 241;
// bram[59647] = 250;
// bram[59648] = 253;
// bram[59649] = 252;
// bram[59650] = 245;
// bram[59651] = 233;
// bram[59652] = 216;
// bram[59653] = 196;
// bram[59654] = 173;
// bram[59655] = 148;
// bram[59656] = 122;
// bram[59657] = 96;
// bram[59658] = 72;
// bram[59659] = 50;
// bram[59660] = 31;
// bram[59661] = 16;
// bram[59662] = 5;
// bram[59663] = 0;
// bram[59664] = 0;
// bram[59665] = 6;
// bram[59666] = 16;
// bram[59667] = 31;
// bram[59668] = 50;
// bram[59669] = 73;
// bram[59670] = 97;
// bram[59671] = 123;
// bram[59672] = 149;
// bram[59673] = 174;
// bram[59674] = 197;
// bram[59675] = 217;
// bram[59676] = 233;
// bram[59677] = 245;
// bram[59678] = 252;
// bram[59679] = 253;
// bram[59680] = 250;
// bram[59681] = 240;
// bram[59682] = 227;
// bram[59683] = 209;
// bram[59684] = 187;
// bram[59685] = 163;
// bram[59686] = 138;
// bram[59687] = 112;
// bram[59688] = 86;
// bram[59689] = 62;
// bram[59690] = 41;
// bram[59691] = 24;
// bram[59692] = 11;
// bram[59693] = 3;
// bram[59694] = 0;
// bram[59695] = 2;
// bram[59696] = 9;
// bram[59697] = 22;
// bram[59698] = 39;
// bram[59699] = 59;
// bram[59700] = 83;
// bram[59701] = 108;
// bram[59702] = 134;
// bram[59703] = 159;
// bram[59704] = 184;
// bram[59705] = 206;
// bram[59706] = 224;
// bram[59707] = 239;
// bram[59708] = 249;
// bram[59709] = 253;
// bram[59710] = 252;
// bram[59711] = 246;
// bram[59712] = 235;
// bram[59713] = 220;
// bram[59714] = 200;
// bram[59715] = 178;
// bram[59716] = 153;
// bram[59717] = 127;
// bram[59718] = 101;
// bram[59719] = 76;
// bram[59720] = 53;
// bram[59721] = 34;
// bram[59722] = 18;
// bram[59723] = 7;
// bram[59724] = 1;
// bram[59725] = 0;
// bram[59726] = 4;
// bram[59727] = 14;
// bram[59728] = 28;
// bram[59729] = 47;
// bram[59730] = 68;
// bram[59731] = 93;
// bram[59732] = 118;
// bram[59733] = 144;
// bram[59734] = 170;
// bram[59735] = 193;
// bram[59736] = 214;
// bram[59737] = 231;
// bram[59738] = 243;
// bram[59739] = 251;
// bram[59740] = 253;
// bram[59741] = 251;
// bram[59742] = 243;
// bram[59743] = 230;
// bram[59744] = 212;
// bram[59745] = 191;
// bram[59746] = 168;
// bram[59747] = 142;
// bram[59748] = 116;
// bram[59749] = 91;
// bram[59750] = 67;
// bram[59751] = 45;
// bram[59752] = 27;
// bram[59753] = 13;
// bram[59754] = 4;
// bram[59755] = 0;
// bram[59756] = 1;
// bram[59757] = 8;
// bram[59758] = 19;
// bram[59759] = 35;
// bram[59760] = 55;
// bram[59761] = 78;
// bram[59762] = 103;
// bram[59763] = 129;
// bram[59764] = 155;
// bram[59765] = 179;
// bram[59766] = 202;
// bram[59767] = 221;
// bram[59768] = 236;
// bram[59769] = 247;
// bram[59770] = 253;
// bram[59771] = 253;
// bram[59772] = 248;
// bram[59773] = 238;
// bram[59774] = 223;
// bram[59775] = 204;
// bram[59776] = 182;
// bram[59777] = 158;
// bram[59778] = 132;
// bram[59779] = 106;
// bram[59780] = 81;
// bram[59781] = 57;
// bram[59782] = 37;
// bram[59783] = 21;
// bram[59784] = 9;
// bram[59785] = 1;
// bram[59786] = 0;
// bram[59787] = 3;
// bram[59788] = 12;
// bram[59789] = 25;
// bram[59790] = 43;
// bram[59791] = 64;
// bram[59792] = 88;
// bram[59793] = 114;
// bram[59794] = 140;
// bram[59795] = 165;
// bram[59796] = 189;
// bram[59797] = 210;
// bram[59798] = 228;
// bram[59799] = 241;
// bram[59800] = 250;
// bram[59801] = 253;
// bram[59802] = 252;
// bram[59803] = 244;
// bram[59804] = 232;
// bram[59805] = 216;
// bram[59806] = 195;
// bram[59807] = 172;
// bram[59808] = 147;
// bram[59809] = 121;
// bram[59810] = 95;
// bram[59811] = 71;
// bram[59812] = 49;
// bram[59813] = 30;
// bram[59814] = 15;
// bram[59815] = 5;
// bram[59816] = 0;
// bram[59817] = 0;
// bram[59818] = 6;
// bram[59819] = 17;
// bram[59820] = 32;
// bram[59821] = 51;
// bram[59822] = 74;
// bram[59823] = 98;
// bram[59824] = 124;
// bram[59825] = 150;
// bram[59826] = 175;
// bram[59827] = 198;
// bram[59828] = 218;
// bram[59829] = 234;
// bram[59830] = 245;
// bram[59831] = 252;
// bram[59832] = 253;
// bram[59833] = 249;
// bram[59834] = 240;
// bram[59835] = 226;
// bram[59836] = 208;
// bram[59837] = 186;
// bram[59838] = 162;
// bram[59839] = 137;
// bram[59840] = 111;
// bram[59841] = 85;
// bram[59842] = 62;
// bram[59843] = 41;
// bram[59844] = 23;
// bram[59845] = 10;
// bram[59846] = 2;
// bram[59847] = 0;
// bram[59848] = 2;
// bram[59849] = 10;
// bram[59850] = 22;
// bram[59851] = 39;
// bram[59852] = 60;
// bram[59853] = 83;
// bram[59854] = 109;
// bram[59855] = 135;
// bram[59856] = 160;
// bram[59857] = 185;
// bram[59858] = 206;
// bram[59859] = 225;
// bram[59860] = 239;
// bram[59861] = 249;
// bram[59862] = 253;
// bram[59863] = 252;
// bram[59864] = 246;
// bram[59865] = 235;
// bram[59866] = 219;
// bram[59867] = 199;
// bram[59868] = 177;
// bram[59869] = 152;
// bram[59870] = 126;
// bram[59871] = 100;
// bram[59872] = 75;
// bram[59873] = 53;
// bram[59874] = 33;
// bram[59875] = 18;
// bram[59876] = 7;
// bram[59877] = 1;
// bram[59878] = 0;
// bram[59879] = 5;
// bram[59880] = 14;
// bram[59881] = 29;
// bram[59882] = 47;
// bram[59883] = 69;
// bram[59884] = 94;
// bram[59885] = 119;
// bram[59886] = 145;
// bram[59887] = 171;
// bram[59888] = 194;
// bram[59889] = 214;
// bram[59890] = 231;
// bram[59891] = 244;
// bram[59892] = 251;
// bram[59893] = 253;
// bram[59894] = 250;
// bram[59895] = 242;
// bram[59896] = 229;
// bram[59897] = 212;
// bram[59898] = 191;
// bram[59899] = 167;
// bram[59900] = 141;
// bram[59901] = 115;
// bram[59902] = 90;
// bram[59903] = 66;
// bram[59904] = 44;
// bram[59905] = 26;
// bram[59906] = 12;
// bram[59907] = 3;
// bram[59908] = 0;
// bram[59909] = 1;
// bram[59910] = 8;
// bram[59911] = 20;
// bram[59912] = 36;
// bram[59913] = 56;
// bram[59914] = 79;
// bram[59915] = 104;
// bram[59916] = 130;
// bram[59917] = 156;
// bram[59918] = 180;
// bram[59919] = 203;
// bram[59920] = 222;
// bram[59921] = 237;
// bram[59922] = 247;
// bram[59923] = 253;
// bram[59924] = 253;
// bram[59925] = 248;
// bram[59926] = 237;
// bram[59927] = 222;
// bram[59928] = 203;
// bram[59929] = 181;
// bram[59930] = 157;
// bram[59931] = 131;
// bram[59932] = 105;
// bram[59933] = 80;
// bram[59934] = 57;
// bram[59935] = 37;
// bram[59936] = 20;
// bram[59937] = 8;
// bram[59938] = 1;
// bram[59939] = 0;
// bram[59940] = 3;
// bram[59941] = 12;
// bram[59942] = 26;
// bram[59943] = 44;
// bram[59944] = 65;
// bram[59945] = 89;
// bram[59946] = 114;
// bram[59947] = 140;
// bram[59948] = 166;
// bram[59949] = 190;
// bram[59950] = 211;
// bram[59951] = 228;
// bram[59952] = 242;
// bram[59953] = 250;
// bram[59954] = 253;
// bram[59955] = 251;
// bram[59956] = 244;
// bram[59957] = 232;
// bram[59958] = 215;
// bram[59959] = 195;
// bram[59960] = 171;
// bram[59961] = 146;
// bram[59962] = 120;
// bram[59963] = 94;
// bram[59964] = 70;
// bram[59965] = 48;
// bram[59966] = 29;
// bram[59967] = 15;
// bram[59968] = 5;
// bram[59969] = 0;
// bram[59970] = 0;
// bram[59971] = 6;
// bram[59972] = 17;
// bram[59973] = 33;
// bram[59974] = 52;
// bram[59975] = 74;
// bram[59976] = 99;
// bram[59977] = 125;
// bram[59978] = 151;
// bram[59979] = 176;
// bram[59980] = 199;
// bram[59981] = 218;
// bram[59982] = 234;
// bram[59983] = 246;
// bram[59984] = 252;
// bram[59985] = 253;
// bram[59986] = 249;
// bram[59987] = 240;
// bram[59988] = 225;
// bram[59989] = 207;
// bram[59990] = 185;
// bram[59991] = 161;
// bram[59992] = 136;
// bram[59993] = 110;
// bram[59994] = 84;
// bram[59995] = 61;
// bram[59996] = 40;
// bram[59997] = 23;
// bram[59998] = 10;
// bram[59999] = 2;
// bram[60000] = 0;
// bram[60001] = 2;
// bram[60002] = 10;
// bram[60003] = 23;
// bram[60004] = 40;
// bram[60005] = 61;
// bram[60006] = 84;
// bram[60007] = 110;
// bram[60008] = 136;
// bram[60009] = 161;
// bram[60010] = 185;
// bram[60011] = 207;
// bram[60012] = 225;
// bram[60013] = 240;
// bram[60014] = 249;
// bram[60015] = 253;
// bram[60016] = 252;
// bram[60017] = 246;
// bram[60018] = 234;
// bram[60019] = 218;
// bram[60020] = 199;
// bram[60021] = 176;
// bram[60022] = 151;
// bram[60023] = 125;
// bram[60024] = 99;
// bram[60025] = 74;
// bram[60026] = 52;
// bram[60027] = 33;
// bram[60028] = 17;
// bram[60029] = 6;
// bram[60030] = 0;
// bram[60031] = 0;
// bram[60032] = 5;
// bram[60033] = 15;
// bram[60034] = 29;
// bram[60035] = 48;
// bram[60036] = 70;
// bram[60037] = 94;
// bram[60038] = 120;
// bram[60039] = 146;
// bram[60040] = 171;
// bram[60041] = 195;
// bram[60042] = 215;
// bram[60043] = 232;
// bram[60044] = 244;
// bram[60045] = 251;
// bram[60046] = 253;
// bram[60047] = 250;
// bram[60048] = 242;
// bram[60049] = 228;
// bram[60050] = 211;
// bram[60051] = 190;
// bram[60052] = 166;
// bram[60053] = 140;
// bram[60054] = 114;
// bram[60055] = 89;
// bram[60056] = 65;
// bram[60057] = 44;
// bram[60058] = 26;
// bram[60059] = 12;
// bram[60060] = 3;
// bram[60061] = 0;
// bram[60062] = 1;
// bram[60063] = 8;
// bram[60064] = 20;
// bram[60065] = 37;
// bram[60066] = 57;
// bram[60067] = 80;
// bram[60068] = 105;
// bram[60069] = 131;
// bram[60070] = 157;
// bram[60071] = 181;
// bram[60072] = 203;
// bram[60073] = 222;
// bram[60074] = 237;
// bram[60075] = 248;
// bram[60076] = 253;
// bram[60077] = 253;
// bram[60078] = 247;
// bram[60079] = 237;
// bram[60080] = 222;
// bram[60081] = 203;
// bram[60082] = 180;
// bram[60083] = 156;
// bram[60084] = 130;
// bram[60085] = 104;
// bram[60086] = 79;
// bram[60087] = 56;
// bram[60088] = 36;
// bram[60089] = 20;
// bram[60090] = 8;
// bram[60091] = 1;
// bram[60092] = 0;
// bram[60093] = 3;
// bram[60094] = 12;
// bram[60095] = 26;
// bram[60096] = 44;
// bram[60097] = 66;
// bram[60098] = 90;
// bram[60099] = 115;
// bram[60100] = 141;
// bram[60101] = 167;
// bram[60102] = 191;
// bram[60103] = 212;
// bram[60104] = 229;
// bram[60105] = 242;
// bram[60106] = 250;
// bram[60107] = 253;
// bram[60108] = 251;
// bram[60109] = 244;
// bram[60110] = 231;
// bram[60111] = 214;
// bram[60112] = 194;
// bram[60113] = 171;
// bram[60114] = 145;
// bram[60115] = 119;
// bram[60116] = 94;
// bram[60117] = 69;
// bram[60118] = 47;
// bram[60119] = 29;
// bram[60120] = 14;
// bram[60121] = 5;
// bram[60122] = 0;
// bram[60123] = 1;
// bram[60124] = 7;
// bram[60125] = 18;
// bram[60126] = 33;
// bram[60127] = 53;
// bram[60128] = 75;
// bram[60129] = 100;
// bram[60130] = 126;
// bram[60131] = 152;
// bram[60132] = 177;
// bram[60133] = 199;
// bram[60134] = 219;
// bram[60135] = 235;
// bram[60136] = 246;
// bram[60137] = 252;
// bram[60138] = 253;
// bram[60139] = 249;
// bram[60140] = 239;
// bram[60141] = 225;
// bram[60142] = 206;
// bram[60143] = 185;
// bram[60144] = 160;
// bram[60145] = 135;
// bram[60146] = 109;
// bram[60147] = 83;
// bram[60148] = 60;
// bram[60149] = 39;
// bram[60150] = 22;
// bram[60151] = 10;
// bram[60152] = 2;
// bram[60153] = 0;
// bram[60154] = 2;
// bram[60155] = 10;
// bram[60156] = 23;
// bram[60157] = 41;
// bram[60158] = 62;
// bram[60159] = 85;
// bram[60160] = 111;
// bram[60161] = 137;
// bram[60162] = 162;
// bram[60163] = 186;
// bram[60164] = 208;
// bram[60165] = 226;
// bram[60166] = 240;
// bram[60167] = 249;
// bram[60168] = 253;
// bram[60169] = 252;
// bram[60170] = 245;
// bram[60171] = 234;
// bram[60172] = 218;
// bram[60173] = 198;
// bram[60174] = 175;
// bram[60175] = 150;
// bram[60176] = 124;
// bram[60177] = 98;
// bram[60178] = 74;
// bram[60179] = 51;
// bram[60180] = 32;
// bram[60181] = 17;
// bram[60182] = 6;
// bram[60183] = 0;
// bram[60184] = 0;
// bram[60185] = 5;
// bram[60186] = 15;
// bram[60187] = 30;
// bram[60188] = 49;
// bram[60189] = 71;
// bram[60190] = 95;
// bram[60191] = 121;
// bram[60192] = 147;
// bram[60193] = 172;
// bram[60194] = 195;
// bram[60195] = 216;
// bram[60196] = 232;
// bram[60197] = 244;
// bram[60198] = 252;
// bram[60199] = 253;
// bram[60200] = 250;
// bram[60201] = 241;
// bram[60202] = 228;
// bram[60203] = 210;
// bram[60204] = 189;
// bram[60205] = 165;
// bram[60206] = 140;
// bram[60207] = 114;
// bram[60208] = 88;
// bram[60209] = 64;
// bram[60210] = 43;
// bram[60211] = 25;
// bram[60212] = 12;
// bram[60213] = 3;
// bram[60214] = 0;
// bram[60215] = 1;
// bram[60216] = 9;
// bram[60217] = 21;
// bram[60218] = 37;
// bram[60219] = 57;
// bram[60220] = 81;
// bram[60221] = 106;
// bram[60222] = 132;
// bram[60223] = 158;
// bram[60224] = 182;
// bram[60225] = 204;
// bram[60226] = 223;
// bram[60227] = 238;
// bram[60228] = 248;
// bram[60229] = 253;
// bram[60230] = 253;
// bram[60231] = 247;
// bram[60232] = 236;
// bram[60233] = 221;
// bram[60234] = 202;
// bram[60235] = 179;
// bram[60236] = 155;
// bram[60237] = 129;
// bram[60238] = 103;
// bram[60239] = 78;
// bram[60240] = 55;
// bram[60241] = 35;
// bram[60242] = 19;
// bram[60243] = 8;
// bram[60244] = 1;
// bram[60245] = 0;
// bram[60246] = 4;
// bram[60247] = 13;
// bram[60248] = 27;
// bram[60249] = 45;
// bram[60250] = 67;
// bram[60251] = 91;
// bram[60252] = 116;
// bram[60253] = 142;
// bram[60254] = 168;
// bram[60255] = 191;
// bram[60256] = 212;
// bram[60257] = 230;
// bram[60258] = 243;
// bram[60259] = 251;
// bram[60260] = 253;
// bram[60261] = 251;
// bram[60262] = 243;
// bram[60263] = 231;
// bram[60264] = 214;
// bram[60265] = 193;
// bram[60266] = 170;
// bram[60267] = 144;
// bram[60268] = 118;
// bram[60269] = 93;
// bram[60270] = 68;
// bram[60271] = 47;
// bram[60272] = 28;
// bram[60273] = 14;
// bram[60274] = 4;
// bram[60275] = 0;
// bram[60276] = 1;
// bram[60277] = 7;
// bram[60278] = 18;
// bram[60279] = 34;
// bram[60280] = 53;
// bram[60281] = 76;
// bram[60282] = 101;
// bram[60283] = 127;
// bram[60284] = 153;
// bram[60285] = 178;
// bram[60286] = 200;
// bram[60287] = 220;
// bram[60288] = 235;
// bram[60289] = 246;
// bram[60290] = 252;
// bram[60291] = 253;
// bram[60292] = 249;
// bram[60293] = 239;
// bram[60294] = 224;
// bram[60295] = 206;
// bram[60296] = 184;
// bram[60297] = 159;
// bram[60298] = 134;
// bram[60299] = 108;
// bram[60300] = 83;
// bram[60301] = 59;
// bram[60302] = 39;
// bram[60303] = 22;
// bram[60304] = 9;
// bram[60305] = 2;
// bram[60306] = 0;
// bram[60307] = 3;
// bram[60308] = 11;
// bram[60309] = 24;
// bram[60310] = 41;
// bram[60311] = 62;
// bram[60312] = 86;
// bram[60313] = 112;
// bram[60314] = 138;
// bram[60315] = 163;
// bram[60316] = 187;
// bram[60317] = 209;
// bram[60318] = 227;
// bram[60319] = 240;
// bram[60320] = 250;
// bram[60321] = 253;
// bram[60322] = 252;
// bram[60323] = 245;
// bram[60324] = 233;
// bram[60325] = 217;
// bram[60326] = 197;
// bram[60327] = 174;
// bram[60328] = 149;
// bram[60329] = 123;
// bram[60330] = 97;
// bram[60331] = 73;
// bram[60332] = 50;
// bram[60333] = 31;
// bram[60334] = 16;
// bram[60335] = 6;
// bram[60336] = 0;
// bram[60337] = 0;
// bram[60338] = 5;
// bram[60339] = 16;
// bram[60340] = 31;
// bram[60341] = 50;
// bram[60342] = 72;
// bram[60343] = 96;
// bram[60344] = 122;
// bram[60345] = 148;
// bram[60346] = 173;
// bram[60347] = 196;
// bram[60348] = 216;
// bram[60349] = 233;
// bram[60350] = 245;
// bram[60351] = 252;
// bram[60352] = 253;
// bram[60353] = 250;
// bram[60354] = 241;
// bram[60355] = 227;
// bram[60356] = 209;
// bram[60357] = 188;
// bram[60358] = 164;
// bram[60359] = 139;
// bram[60360] = 113;
// bram[60361] = 87;
// bram[60362] = 63;
// bram[60363] = 42;
// bram[60364] = 25;
// bram[60365] = 11;
// bram[60366] = 3;
// bram[60367] = 0;
// bram[60368] = 2;
// bram[60369] = 9;
// bram[60370] = 21;
// bram[60371] = 38;
// bram[60372] = 58;
// bram[60373] = 82;
// bram[60374] = 107;
// bram[60375] = 133;
// bram[60376] = 158;
// bram[60377] = 183;
// bram[60378] = 205;
// bram[60379] = 224;
// bram[60380] = 238;
// bram[60381] = 248;
// bram[60382] = 253;
// bram[60383] = 253;
// bram[60384] = 247;
// bram[60385] = 236;
// bram[60386] = 221;
// bram[60387] = 201;
// bram[60388] = 179;
// bram[60389] = 154;
// bram[60390] = 128;
// bram[60391] = 102;
// bram[60392] = 77;
// bram[60393] = 54;
// bram[60394] = 35;
// bram[60395] = 19;
// bram[60396] = 7;
// bram[60397] = 1;
// bram[60398] = 0;
// bram[60399] = 4;
// bram[60400] = 13;
// bram[60401] = 27;
// bram[60402] = 46;
// bram[60403] = 67;
// bram[60404] = 92;
// bram[60405] = 117;
// bram[60406] = 143;
// bram[60407] = 169;
// bram[60408] = 192;
// bram[60409] = 213;
// bram[60410] = 230;
// bram[60411] = 243;
// bram[60412] = 251;
// bram[60413] = 253;
// bram[60414] = 251;
// bram[60415] = 243;
// bram[60416] = 230;
// bram[60417] = 213;
// bram[60418] = 192;
// bram[60419] = 169;
// bram[60420] = 143;
// bram[60421] = 117;
// bram[60422] = 92;
// bram[60423] = 68;
// bram[60424] = 46;
// bram[60425] = 28;
// bram[60426] = 13;
// bram[60427] = 4;
// bram[60428] = 0;
// bram[60429] = 1;
// bram[60430] = 7;
// bram[60431] = 19;
// bram[60432] = 34;
// bram[60433] = 54;
// bram[60434] = 77;
// bram[60435] = 102;
// bram[60436] = 128;
// bram[60437] = 154;
// bram[60438] = 178;
// bram[60439] = 201;
// bram[60440] = 220;
// bram[60441] = 236;
// bram[60442] = 247;
// bram[60443] = 253;
// bram[60444] = 253;
// bram[60445] = 248;
// bram[60446] = 238;
// bram[60447] = 224;
// bram[60448] = 205;
// bram[60449] = 183;
// bram[60450] = 159;
// bram[60451] = 133;
// bram[60452] = 107;
// bram[60453] = 82;
// bram[60454] = 58;
// bram[60455] = 38;
// bram[60456] = 21;
// bram[60457] = 9;
// bram[60458] = 2;
// bram[60459] = 0;
// bram[60460] = 3;
// bram[60461] = 11;
// bram[60462] = 25;
// bram[60463] = 42;
// bram[60464] = 63;
// bram[60465] = 87;
// bram[60466] = 112;
// bram[60467] = 139;
// bram[60468] = 164;
// bram[60469] = 188;
// bram[60470] = 209;
// bram[60471] = 227;
// bram[60472] = 241;
// bram[60473] = 250;
// bram[60474] = 253;
// bram[60475] = 252;
// bram[60476] = 245;
// bram[60477] = 233;
// bram[60478] = 217;
// bram[60479] = 196;
// bram[60480] = 173;
// bram[60481] = 148;
// bram[60482] = 122;
// bram[60483] = 96;
// bram[60484] = 72;
// bram[60485] = 50;
// bram[60486] = 31;
// bram[60487] = 16;
// bram[60488] = 5;
// bram[60489] = 0;
// bram[60490] = 0;
// bram[60491] = 6;
// bram[60492] = 16;
// bram[60493] = 31;
// bram[60494] = 50;
// bram[60495] = 73;
// bram[60496] = 97;
// bram[60497] = 123;
// bram[60498] = 149;
// bram[60499] = 174;
// bram[60500] = 197;
// bram[60501] = 217;
// bram[60502] = 233;
// bram[60503] = 245;
// bram[60504] = 252;
// bram[60505] = 253;
// bram[60506] = 250;
// bram[60507] = 241;
// bram[60508] = 227;
// bram[60509] = 209;
// bram[60510] = 187;
// bram[60511] = 163;
// bram[60512] = 138;
// bram[60513] = 112;
// bram[60514] = 86;
// bram[60515] = 62;
// bram[60516] = 41;
// bram[60517] = 24;
// bram[60518] = 11;
// bram[60519] = 3;
// bram[60520] = 0;
// bram[60521] = 2;
// bram[60522] = 9;
// bram[60523] = 22;
// bram[60524] = 39;
// bram[60525] = 59;
// bram[60526] = 82;
// bram[60527] = 108;
// bram[60528] = 134;
// bram[60529] = 159;
// bram[60530] = 184;
// bram[60531] = 206;
// bram[60532] = 224;
// bram[60533] = 239;
// bram[60534] = 248;
// bram[60535] = 253;
// bram[60536] = 252;
// bram[60537] = 246;
// bram[60538] = 235;
// bram[60539] = 220;
// bram[60540] = 200;
// bram[60541] = 178;
// bram[60542] = 153;
// bram[60543] = 127;
// bram[60544] = 101;
// bram[60545] = 76;
// bram[60546] = 54;
// bram[60547] = 34;
// bram[60548] = 18;
// bram[60549] = 7;
// bram[60550] = 1;
// bram[60551] = 0;
// bram[60552] = 4;
// bram[60553] = 14;
// bram[60554] = 28;
// bram[60555] = 47;
// bram[60556] = 68;
// bram[60557] = 93;
// bram[60558] = 118;
// bram[60559] = 144;
// bram[60560] = 170;
// bram[60561] = 193;
// bram[60562] = 214;
// bram[60563] = 231;
// bram[60564] = 243;
// bram[60565] = 251;
// bram[60566] = 253;
// bram[60567] = 251;
// bram[60568] = 243;
// bram[60569] = 230;
// bram[60570] = 212;
// bram[60571] = 191;
// bram[60572] = 168;
// bram[60573] = 142;
// bram[60574] = 116;
// bram[60575] = 91;
// bram[60576] = 67;
// bram[60577] = 45;
// bram[60578] = 27;
// bram[60579] = 13;
// bram[60580] = 4;
// bram[60581] = 0;
// bram[60582] = 1;
// bram[60583] = 8;
// bram[60584] = 19;
// bram[60585] = 35;
// bram[60586] = 55;
// bram[60587] = 78;
// bram[60588] = 103;
// bram[60589] = 129;
// bram[60590] = 155;
// bram[60591] = 179;
// bram[60592] = 202;
// bram[60593] = 221;
// bram[60594] = 236;
// bram[60595] = 247;
// bram[60596] = 253;
// bram[60597] = 253;
// bram[60598] = 248;
// bram[60599] = 238;
// bram[60600] = 223;
// bram[60601] = 204;
// bram[60602] = 182;
// bram[60603] = 158;
// bram[60604] = 132;
// bram[60605] = 106;
// bram[60606] = 81;
// bram[60607] = 58;
// bram[60608] = 37;
// bram[60609] = 21;
// bram[60610] = 9;
// bram[60611] = 1;
// bram[60612] = 0;
// bram[60613] = 3;
// bram[60614] = 12;
// bram[60615] = 25;
// bram[60616] = 43;
// bram[60617] = 64;
// bram[60618] = 88;
// bram[60619] = 113;
// bram[60620] = 139;
// bram[60621] = 165;
// bram[60622] = 189;
// bram[60623] = 210;
// bram[60624] = 228;
// bram[60625] = 241;
// bram[60626] = 250;
// bram[60627] = 253;
// bram[60628] = 252;
// bram[60629] = 244;
// bram[60630] = 232;
// bram[60631] = 216;
// bram[60632] = 196;
// bram[60633] = 172;
// bram[60634] = 147;
// bram[60635] = 121;
// bram[60636] = 95;
// bram[60637] = 71;
// bram[60638] = 49;
// bram[60639] = 30;
// bram[60640] = 15;
// bram[60641] = 5;
// bram[60642] = 0;
// bram[60643] = 0;
// bram[60644] = 6;
// bram[60645] = 17;
// bram[60646] = 32;
// bram[60647] = 51;
// bram[60648] = 74;
// bram[60649] = 98;
// bram[60650] = 124;
// bram[60651] = 150;
// bram[60652] = 175;
// bram[60653] = 198;
// bram[60654] = 218;
// bram[60655] = 234;
// bram[60656] = 245;
// bram[60657] = 252;
// bram[60658] = 253;
// bram[60659] = 249;
// bram[60660] = 240;
// bram[60661] = 226;
// bram[60662] = 208;
// bram[60663] = 186;
// bram[60664] = 162;
// bram[60665] = 137;
// bram[60666] = 111;
// bram[60667] = 85;
// bram[60668] = 62;
// bram[60669] = 41;
// bram[60670] = 23;
// bram[60671] = 10;
// bram[60672] = 2;
// bram[60673] = 0;
// bram[60674] = 2;
// bram[60675] = 10;
// bram[60676] = 22;
// bram[60677] = 39;
// bram[60678] = 60;
// bram[60679] = 83;
// bram[60680] = 109;
// bram[60681] = 135;
// bram[60682] = 160;
// bram[60683] = 185;
// bram[60684] = 206;
// bram[60685] = 225;
// bram[60686] = 239;
// bram[60687] = 249;
// bram[60688] = 253;
// bram[60689] = 252;
// bram[60690] = 246;
// bram[60691] = 235;
// bram[60692] = 219;
// bram[60693] = 200;
// bram[60694] = 177;
// bram[60695] = 152;
// bram[60696] = 126;
// bram[60697] = 100;
// bram[60698] = 75;
// bram[60699] = 53;
// bram[60700] = 33;
// bram[60701] = 18;
// bram[60702] = 7;
// bram[60703] = 1;
// bram[60704] = 0;
// bram[60705] = 4;
// bram[60706] = 14;
// bram[60707] = 29;
// bram[60708] = 47;
// bram[60709] = 69;
// bram[60710] = 93;
// bram[60711] = 119;
// bram[60712] = 145;
// bram[60713] = 170;
// bram[60714] = 194;
// bram[60715] = 214;
// bram[60716] = 231;
// bram[60717] = 244;
// bram[60718] = 251;
// bram[60719] = 253;
// bram[60720] = 250;
// bram[60721] = 242;
// bram[60722] = 229;
// bram[60723] = 212;
// bram[60724] = 191;
// bram[60725] = 167;
// bram[60726] = 142;
// bram[60727] = 115;
// bram[60728] = 90;
// bram[60729] = 66;
// bram[60730] = 44;
// bram[60731] = 26;
// bram[60732] = 13;
// bram[60733] = 4;
// bram[60734] = 0;
// bram[60735] = 1;
// bram[60736] = 8;
// bram[60737] = 20;
// bram[60738] = 36;
// bram[60739] = 56;
// bram[60740] = 79;
// bram[60741] = 104;
// bram[60742] = 130;
// bram[60743] = 156;
// bram[60744] = 180;
// bram[60745] = 203;
// bram[60746] = 222;
// bram[60747] = 237;
// bram[60748] = 247;
// bram[60749] = 253;
// bram[60750] = 253;
// bram[60751] = 248;
// bram[60752] = 237;
// bram[60753] = 222;
// bram[60754] = 203;
// bram[60755] = 181;
// bram[60756] = 157;
// bram[60757] = 131;
// bram[60758] = 105;
// bram[60759] = 80;
// bram[60760] = 57;
// bram[60761] = 37;
// bram[60762] = 20;
// bram[60763] = 8;
// bram[60764] = 1;
// bram[60765] = 0;
// bram[60766] = 3;
// bram[60767] = 12;
// bram[60768] = 26;
// bram[60769] = 44;
// bram[60770] = 65;
// bram[60771] = 89;
// bram[60772] = 114;
// bram[60773] = 140;
// bram[60774] = 166;
// bram[60775] = 190;
// bram[60776] = 211;
// bram[60777] = 228;
// bram[60778] = 242;
// bram[60779] = 250;
// bram[60780] = 253;
// bram[60781] = 251;
// bram[60782] = 244;
// bram[60783] = 232;
// bram[60784] = 215;
// bram[60785] = 195;
// bram[60786] = 171;
// bram[60787] = 146;
// bram[60788] = 120;
// bram[60789] = 95;
// bram[60790] = 70;
// bram[60791] = 48;
// bram[60792] = 29;
// bram[60793] = 15;
// bram[60794] = 5;
// bram[60795] = 0;
// bram[60796] = 0;
// bram[60797] = 6;
// bram[60798] = 17;
// bram[60799] = 32;
// bram[60800] = 52;
// bram[60801] = 74;
// bram[60802] = 99;
// bram[60803] = 125;
// bram[60804] = 151;
// bram[60805] = 176;
// bram[60806] = 199;
// bram[60807] = 218;
// bram[60808] = 234;
// bram[60809] = 246;
// bram[60810] = 252;
// bram[60811] = 253;
// bram[60812] = 249;
// bram[60813] = 240;
// bram[60814] = 226;
// bram[60815] = 207;
// bram[60816] = 186;
// bram[60817] = 161;
// bram[60818] = 136;
// bram[60819] = 110;
// bram[60820] = 84;
// bram[60821] = 61;
// bram[60822] = 40;
// bram[60823] = 23;
// bram[60824] = 10;
// bram[60825] = 2;
// bram[60826] = 0;
// bram[60827] = 2;
// bram[60828] = 10;
// bram[60829] = 23;
// bram[60830] = 40;
// bram[60831] = 61;
// bram[60832] = 84;
// bram[60833] = 110;
// bram[60834] = 136;
// bram[60835] = 161;
// bram[60836] = 185;
// bram[60837] = 207;
// bram[60838] = 225;
// bram[60839] = 240;
// bram[60840] = 249;
// bram[60841] = 253;
// bram[60842] = 252;
// bram[60843] = 246;
// bram[60844] = 234;
// bram[60845] = 219;
// bram[60846] = 199;
// bram[60847] = 176;
// bram[60848] = 151;
// bram[60849] = 125;
// bram[60850] = 99;
// bram[60851] = 75;
// bram[60852] = 52;
// bram[60853] = 33;
// bram[60854] = 17;
// bram[60855] = 6;
// bram[60856] = 0;
// bram[60857] = 0;
// bram[60858] = 5;
// bram[60859] = 15;
// bram[60860] = 29;
// bram[60861] = 48;
// bram[60862] = 70;
// bram[60863] = 94;
// bram[60864] = 120;
// bram[60865] = 146;
// bram[60866] = 171;
// bram[60867] = 195;
// bram[60868] = 215;
// bram[60869] = 232;
// bram[60870] = 244;
// bram[60871] = 251;
// bram[60872] = 253;
// bram[60873] = 250;
// bram[60874] = 242;
// bram[60875] = 229;
// bram[60876] = 211;
// bram[60877] = 190;
// bram[60878] = 166;
// bram[60879] = 141;
// bram[60880] = 115;
// bram[60881] = 89;
// bram[60882] = 65;
// bram[60883] = 44;
// bram[60884] = 26;
// bram[60885] = 12;
// bram[60886] = 3;
// bram[60887] = 0;
// bram[60888] = 1;
// bram[60889] = 8;
// bram[60890] = 20;
// bram[60891] = 36;
// bram[60892] = 57;
// bram[60893] = 80;
// bram[60894] = 105;
// bram[60895] = 131;
// bram[60896] = 157;
// bram[60897] = 181;
// bram[60898] = 203;
// bram[60899] = 222;
// bram[60900] = 237;
// bram[60901] = 248;
// bram[60902] = 253;
// bram[60903] = 253;
// bram[60904] = 247;
// bram[60905] = 237;
// bram[60906] = 222;
// bram[60907] = 203;
// bram[60908] = 180;
// bram[60909] = 156;
// bram[60910] = 130;
// bram[60911] = 104;
// bram[60912] = 79;
// bram[60913] = 56;
// bram[60914] = 36;
// bram[60915] = 20;
// bram[60916] = 8;
// bram[60917] = 1;
// bram[60918] = 0;
// bram[60919] = 3;
// bram[60920] = 12;
// bram[60921] = 26;
// bram[60922] = 44;
// bram[60923] = 66;
// bram[60924] = 90;
// bram[60925] = 115;
// bram[60926] = 141;
// bram[60927] = 167;
// bram[60928] = 190;
// bram[60929] = 211;
// bram[60930] = 229;
// bram[60931] = 242;
// bram[60932] = 250;
// bram[60933] = 253;
// bram[60934] = 251;
// bram[60935] = 244;
// bram[60936] = 231;
// bram[60937] = 214;
// bram[60938] = 194;
// bram[60939] = 171;
// bram[60940] = 145;
// bram[60941] = 119;
// bram[60942] = 94;
// bram[60943] = 69;
// bram[60944] = 47;
// bram[60945] = 29;
// bram[60946] = 14;
// bram[60947] = 5;
// bram[60948] = 0;
// bram[60949] = 1;
// bram[60950] = 7;
// bram[60951] = 18;
// bram[60952] = 33;
// bram[60953] = 53;
// bram[60954] = 75;
// bram[60955] = 100;
// bram[60956] = 126;
// bram[60957] = 152;
// bram[60958] = 177;
// bram[60959] = 199;
// bram[60960] = 219;
// bram[60961] = 235;
// bram[60962] = 246;
// bram[60963] = 252;
// bram[60964] = 253;
// bram[60965] = 249;
// bram[60966] = 239;
// bram[60967] = 225;
// bram[60968] = 207;
// bram[60969] = 185;
// bram[60970] = 160;
// bram[60971] = 135;
// bram[60972] = 109;
// bram[60973] = 84;
// bram[60974] = 60;
// bram[60975] = 39;
// bram[60976] = 22;
// bram[60977] = 10;
// bram[60978] = 2;
// bram[60979] = 0;
// bram[60980] = 2;
// bram[60981] = 10;
// bram[60982] = 23;
// bram[60983] = 41;
// bram[60984] = 62;
// bram[60985] = 85;
// bram[60986] = 110;
// bram[60987] = 137;
// bram[60988] = 162;
// bram[60989] = 186;
// bram[60990] = 208;
// bram[60991] = 226;
// bram[60992] = 240;
// bram[60993] = 249;
// bram[60994] = 253;
// bram[60995] = 252;
// bram[60996] = 246;
// bram[60997] = 234;
// bram[60998] = 218;
// bram[60999] = 198;
// bram[61000] = 175;
// bram[61001] = 150;
// bram[61002] = 124;
// bram[61003] = 98;
// bram[61004] = 74;
// bram[61005] = 51;
// bram[61006] = 32;
// bram[61007] = 17;
// bram[61008] = 6;
// bram[61009] = 0;
// bram[61010] = 0;
// bram[61011] = 5;
// bram[61012] = 15;
// bram[61013] = 30;
// bram[61014] = 49;
// bram[61015] = 71;
// bram[61016] = 95;
// bram[61017] = 121;
// bram[61018] = 147;
// bram[61019] = 172;
// bram[61020] = 195;
// bram[61021] = 216;
// bram[61022] = 232;
// bram[61023] = 244;
// bram[61024] = 252;
// bram[61025] = 253;
// bram[61026] = 250;
// bram[61027] = 241;
// bram[61028] = 228;
// bram[61029] = 210;
// bram[61030] = 189;
// bram[61031] = 165;
// bram[61032] = 140;
// bram[61033] = 114;
// bram[61034] = 88;
// bram[61035] = 64;
// bram[61036] = 43;
// bram[61037] = 25;
// bram[61038] = 12;
// bram[61039] = 3;
// bram[61040] = 0;
// bram[61041] = 1;
// bram[61042] = 9;
// bram[61043] = 21;
// bram[61044] = 37;
// bram[61045] = 57;
// bram[61046] = 81;
// bram[61047] = 106;
// bram[61048] = 132;
// bram[61049] = 157;
// bram[61050] = 182;
// bram[61051] = 204;
// bram[61052] = 223;
// bram[61053] = 238;
// bram[61054] = 248;
// bram[61055] = 253;
// bram[61056] = 253;
// bram[61057] = 247;
// bram[61058] = 236;
// bram[61059] = 221;
// bram[61060] = 202;
// bram[61061] = 180;
// bram[61062] = 155;
// bram[61063] = 129;
// bram[61064] = 103;
// bram[61065] = 78;
// bram[61066] = 55;
// bram[61067] = 35;
// bram[61068] = 19;
// bram[61069] = 8;
// bram[61070] = 1;
// bram[61071] = 0;
// bram[61072] = 4;
// bram[61073] = 13;
// bram[61074] = 27;
// bram[61075] = 45;
// bram[61076] = 67;
// bram[61077] = 91;
// bram[61078] = 116;
// bram[61079] = 142;
// bram[61080] = 168;
// bram[61081] = 191;
// bram[61082] = 212;
// bram[61083] = 230;
// bram[61084] = 242;
// bram[61085] = 251;
// bram[61086] = 253;
// bram[61087] = 251;
// bram[61088] = 243;
// bram[61089] = 231;
// bram[61090] = 214;
// bram[61091] = 193;
// bram[61092] = 170;
// bram[61093] = 144;
// bram[61094] = 118;
// bram[61095] = 93;
// bram[61096] = 68;
// bram[61097] = 47;
// bram[61098] = 28;
// bram[61099] = 14;
// bram[61100] = 4;
// bram[61101] = 0;
// bram[61102] = 1;
// bram[61103] = 7;
// bram[61104] = 18;
// bram[61105] = 34;
// bram[61106] = 53;
// bram[61107] = 76;
// bram[61108] = 101;
// bram[61109] = 127;
// bram[61110] = 153;
// bram[61111] = 178;
// bram[61112] = 200;
// bram[61113] = 220;
// bram[61114] = 235;
// bram[61115] = 246;
// bram[61116] = 252;
// bram[61117] = 253;
// bram[61118] = 249;
// bram[61119] = 239;
// bram[61120] = 224;
// bram[61121] = 206;
// bram[61122] = 184;
// bram[61123] = 160;
// bram[61124] = 134;
// bram[61125] = 108;
// bram[61126] = 83;
// bram[61127] = 59;
// bram[61128] = 39;
// bram[61129] = 22;
// bram[61130] = 9;
// bram[61131] = 2;
// bram[61132] = 0;
// bram[61133] = 3;
// bram[61134] = 11;
// bram[61135] = 24;
// bram[61136] = 41;
// bram[61137] = 62;
// bram[61138] = 86;
// bram[61139] = 111;
// bram[61140] = 137;
// bram[61141] = 163;
// bram[61142] = 187;
// bram[61143] = 209;
// bram[61144] = 227;
// bram[61145] = 240;
// bram[61146] = 249;
// bram[61147] = 253;
// bram[61148] = 252;
// bram[61149] = 245;
// bram[61150] = 233;
// bram[61151] = 217;
// bram[61152] = 197;
// bram[61153] = 174;
// bram[61154] = 149;
// bram[61155] = 123;
// bram[61156] = 97;
// bram[61157] = 73;
// bram[61158] = 50;
// bram[61159] = 31;
// bram[61160] = 16;
// bram[61161] = 6;
// bram[61162] = 0;
// bram[61163] = 0;
// bram[61164] = 5;
// bram[61165] = 16;
// bram[61166] = 31;
// bram[61167] = 49;
// bram[61168] = 72;
// bram[61169] = 96;
// bram[61170] = 122;
// bram[61171] = 148;
// bram[61172] = 173;
// bram[61173] = 196;
// bram[61174] = 216;
// bram[61175] = 233;
// bram[61176] = 245;
// bram[61177] = 252;
// bram[61178] = 253;
// bram[61179] = 250;
// bram[61180] = 241;
// bram[61181] = 227;
// bram[61182] = 210;
// bram[61183] = 188;
// bram[61184] = 164;
// bram[61185] = 139;
// bram[61186] = 113;
// bram[61187] = 87;
// bram[61188] = 63;
// bram[61189] = 42;
// bram[61190] = 25;
// bram[61191] = 11;
// bram[61192] = 3;
// bram[61193] = 0;
// bram[61194] = 2;
// bram[61195] = 9;
// bram[61196] = 21;
// bram[61197] = 38;
// bram[61198] = 58;
// bram[61199] = 81;
// bram[61200] = 107;
// bram[61201] = 133;
// bram[61202] = 158;
// bram[61203] = 183;
// bram[61204] = 205;
// bram[61205] = 224;
// bram[61206] = 238;
// bram[61207] = 248;
// bram[61208] = 253;
// bram[61209] = 253;
// bram[61210] = 247;
// bram[61211] = 236;
// bram[61212] = 221;
// bram[61213] = 201;
// bram[61214] = 179;
// bram[61215] = 154;
// bram[61216] = 128;
// bram[61217] = 102;
// bram[61218] = 77;
// bram[61219] = 54;
// bram[61220] = 35;
// bram[61221] = 19;
// bram[61222] = 7;
// bram[61223] = 1;
// bram[61224] = 0;
// bram[61225] = 4;
// bram[61226] = 13;
// bram[61227] = 27;
// bram[61228] = 46;
// bram[61229] = 67;
// bram[61230] = 92;
// bram[61231] = 117;
// bram[61232] = 143;
// bram[61233] = 169;
// bram[61234] = 192;
// bram[61235] = 213;
// bram[61236] = 230;
// bram[61237] = 243;
// bram[61238] = 251;
// bram[61239] = 253;
// bram[61240] = 251;
// bram[61241] = 243;
// bram[61242] = 230;
// bram[61243] = 213;
// bram[61244] = 192;
// bram[61245] = 169;
// bram[61246] = 144;
// bram[61247] = 117;
// bram[61248] = 92;
// bram[61249] = 68;
// bram[61250] = 46;
// bram[61251] = 28;
// bram[61252] = 13;
// bram[61253] = 4;
// bram[61254] = 0;
// bram[61255] = 1;
// bram[61256] = 7;
// bram[61257] = 19;
// bram[61258] = 34;
// bram[61259] = 54;
// bram[61260] = 77;
// bram[61261] = 102;
// bram[61262] = 128;
// bram[61263] = 154;
// bram[61264] = 178;
// bram[61265] = 201;
// bram[61266] = 220;
// bram[61267] = 236;
// bram[61268] = 247;
// bram[61269] = 253;
// bram[61270] = 253;
// bram[61271] = 248;
// bram[61272] = 238;
// bram[61273] = 224;
// bram[61274] = 205;
// bram[61275] = 183;
// bram[61276] = 159;
// bram[61277] = 133;
// bram[61278] = 107;
// bram[61279] = 82;
// bram[61280] = 58;
// bram[61281] = 38;
// bram[61282] = 21;
// bram[61283] = 9;
// bram[61284] = 2;
// bram[61285] = 0;
// bram[61286] = 3;
// bram[61287] = 11;
// bram[61288] = 24;
// bram[61289] = 42;
// bram[61290] = 63;
// bram[61291] = 87;
// bram[61292] = 112;
// bram[61293] = 138;
// bram[61294] = 164;
// bram[61295] = 188;
// bram[61296] = 209;
// bram[61297] = 227;
// bram[61298] = 241;
// bram[61299] = 250;
// bram[61300] = 253;
// bram[61301] = 252;
// bram[61302] = 245;
// bram[61303] = 233;
// bram[61304] = 217;
// bram[61305] = 196;
// bram[61306] = 173;
// bram[61307] = 148;
// bram[61308] = 122;
// bram[61309] = 97;
// bram[61310] = 72;
// bram[61311] = 50;
// bram[61312] = 31;
// bram[61313] = 16;
// bram[61314] = 5;
// bram[61315] = 0;
// bram[61316] = 0;
// bram[61317] = 6;
// bram[61318] = 16;
// bram[61319] = 31;
// bram[61320] = 50;
// bram[61321] = 73;
// bram[61322] = 97;
// bram[61323] = 123;
// bram[61324] = 149;
// bram[61325] = 174;
// bram[61326] = 197;
// bram[61327] = 217;
// bram[61328] = 233;
// bram[61329] = 245;
// bram[61330] = 252;
// bram[61331] = 253;
// bram[61332] = 250;
// bram[61333] = 241;
// bram[61334] = 227;
// bram[61335] = 209;
// bram[61336] = 187;
// bram[61337] = 163;
// bram[61338] = 138;
// bram[61339] = 112;
// bram[61340] = 86;
// bram[61341] = 63;
// bram[61342] = 42;
// bram[61343] = 24;
// bram[61344] = 11;
// bram[61345] = 3;
// bram[61346] = 0;
// bram[61347] = 2;
// bram[61348] = 9;
// bram[61349] = 22;
// bram[61350] = 38;
// bram[61351] = 59;
// bram[61352] = 82;
// bram[61353] = 108;
// bram[61354] = 134;
// bram[61355] = 159;
// bram[61356] = 184;
// bram[61357] = 206;
// bram[61358] = 224;
// bram[61359] = 239;
// bram[61360] = 248;
// bram[61361] = 253;
// bram[61362] = 252;
// bram[61363] = 247;
// bram[61364] = 236;
// bram[61365] = 220;
// bram[61366] = 200;
// bram[61367] = 178;
// bram[61368] = 153;
// bram[61369] = 127;
// bram[61370] = 101;
// bram[61371] = 76;
// bram[61372] = 54;
// bram[61373] = 34;
// bram[61374] = 18;
// bram[61375] = 7;
// bram[61376] = 1;
// bram[61377] = 0;
// bram[61378] = 4;
// bram[61379] = 14;
// bram[61380] = 28;
// bram[61381] = 46;
// bram[61382] = 68;
// bram[61383] = 92;
// bram[61384] = 118;
// bram[61385] = 144;
// bram[61386] = 169;
// bram[61387] = 193;
// bram[61388] = 214;
// bram[61389] = 231;
// bram[61390] = 243;
// bram[61391] = 251;
// bram[61392] = 253;
// bram[61393] = 251;
// bram[61394] = 243;
// bram[61395] = 230;
// bram[61396] = 212;
// bram[61397] = 192;
// bram[61398] = 168;
// bram[61399] = 143;
// bram[61400] = 117;
// bram[61401] = 91;
// bram[61402] = 67;
// bram[61403] = 45;
// bram[61404] = 27;
// bram[61405] = 13;
// bram[61406] = 4;
// bram[61407] = 0;
// bram[61408] = 1;
// bram[61409] = 7;
// bram[61410] = 19;
// bram[61411] = 35;
// bram[61412] = 55;
// bram[61413] = 78;
// bram[61414] = 103;
// bram[61415] = 129;
// bram[61416] = 155;
// bram[61417] = 179;
// bram[61418] = 202;
// bram[61419] = 221;
// bram[61420] = 236;
// bram[61421] = 247;
// bram[61422] = 253;
// bram[61423] = 253;
// bram[61424] = 248;
// bram[61425] = 238;
// bram[61426] = 223;
// bram[61427] = 204;
// bram[61428] = 182;
// bram[61429] = 158;
// bram[61430] = 132;
// bram[61431] = 106;
// bram[61432] = 81;
// bram[61433] = 58;
// bram[61434] = 37;
// bram[61435] = 21;
// bram[61436] = 9;
// bram[61437] = 1;
// bram[61438] = 0;
// bram[61439] = 3;
// bram[61440] = 12;
// bram[61441] = 25;
// bram[61442] = 43;
// bram[61443] = 64;
// bram[61444] = 88;
// bram[61445] = 113;
// bram[61446] = 139;
// bram[61447] = 165;
// bram[61448] = 189;
// bram[61449] = 210;
// bram[61450] = 228;
// bram[61451] = 241;
// bram[61452] = 250;
// bram[61453] = 253;
// bram[61454] = 252;
// bram[61455] = 244;
// bram[61456] = 232;
// bram[61457] = 216;
// bram[61458] = 196;
// bram[61459] = 172;
// bram[61460] = 147;
// bram[61461] = 121;
// bram[61462] = 96;
// bram[61463] = 71;
// bram[61464] = 49;
// bram[61465] = 30;
// bram[61466] = 15;
// bram[61467] = 5;
// bram[61468] = 0;
// bram[61469] = 0;
// bram[61470] = 6;
// bram[61471] = 17;
// bram[61472] = 32;
// bram[61473] = 51;
// bram[61474] = 73;
// bram[61475] = 98;
// bram[61476] = 124;
// bram[61477] = 150;
// bram[61478] = 175;
// bram[61479] = 198;
// bram[61480] = 218;
// bram[61481] = 234;
// bram[61482] = 245;
// bram[61483] = 252;
// bram[61484] = 253;
// bram[61485] = 249;
// bram[61486] = 240;
// bram[61487] = 226;
// bram[61488] = 208;
// bram[61489] = 186;
// bram[61490] = 162;
// bram[61491] = 137;
// bram[61492] = 111;
// bram[61493] = 85;
// bram[61494] = 62;
// bram[61495] = 41;
// bram[61496] = 24;
// bram[61497] = 11;
// bram[61498] = 2;
// bram[61499] = 0;
// bram[61500] = 2;
// bram[61501] = 10;
// bram[61502] = 22;
// bram[61503] = 39;
// bram[61504] = 60;
// bram[61505] = 83;
// bram[61506] = 109;
// bram[61507] = 135;
// bram[61508] = 160;
// bram[61509] = 184;
// bram[61510] = 206;
// bram[61511] = 225;
// bram[61512] = 239;
// bram[61513] = 249;
// bram[61514] = 253;
// bram[61515] = 252;
// bram[61516] = 246;
// bram[61517] = 235;
// bram[61518] = 219;
// bram[61519] = 200;
// bram[61520] = 177;
// bram[61521] = 152;
// bram[61522] = 126;
// bram[61523] = 100;
// bram[61524] = 76;
// bram[61525] = 53;
// bram[61526] = 33;
// bram[61527] = 18;
// bram[61528] = 7;
// bram[61529] = 1;
// bram[61530] = 0;
// bram[61531] = 4;
// bram[61532] = 14;
// bram[61533] = 29;
// bram[61534] = 47;
// bram[61535] = 69;
// bram[61536] = 93;
// bram[61537] = 119;
// bram[61538] = 145;
// bram[61539] = 170;
// bram[61540] = 194;
// bram[61541] = 214;
// bram[61542] = 231;
// bram[61543] = 244;
// bram[61544] = 251;
// bram[61545] = 253;
// bram[61546] = 250;
// bram[61547] = 242;
// bram[61548] = 229;
// bram[61549] = 212;
// bram[61550] = 191;
// bram[61551] = 167;
// bram[61552] = 142;
// bram[61553] = 116;
// bram[61554] = 90;
// bram[61555] = 66;
// bram[61556] = 44;
// bram[61557] = 26;
// bram[61558] = 13;
// bram[61559] = 4;
// bram[61560] = 0;
// bram[61561] = 1;
// bram[61562] = 8;
// bram[61563] = 20;
// bram[61564] = 36;
// bram[61565] = 56;
// bram[61566] = 79;
// bram[61567] = 104;
// bram[61568] = 130;
// bram[61569] = 156;
// bram[61570] = 180;
// bram[61571] = 202;
// bram[61572] = 222;
// bram[61573] = 237;
// bram[61574] = 247;
// bram[61575] = 253;
// bram[61576] = 253;
// bram[61577] = 248;
// bram[61578] = 237;
// bram[61579] = 223;
// bram[61580] = 204;
// bram[61581] = 181;
// bram[61582] = 157;
// bram[61583] = 131;
// bram[61584] = 105;
// bram[61585] = 80;
// bram[61586] = 57;
// bram[61587] = 37;
// bram[61588] = 20;
// bram[61589] = 8;
// bram[61590] = 1;
// bram[61591] = 0;
// bram[61592] = 3;
// bram[61593] = 12;
// bram[61594] = 26;
// bram[61595] = 43;
// bram[61596] = 65;
// bram[61597] = 89;
// bram[61598] = 114;
// bram[61599] = 140;
// bram[61600] = 166;
// bram[61601] = 190;
// bram[61602] = 211;
// bram[61603] = 228;
// bram[61604] = 242;
// bram[61605] = 250;
// bram[61606] = 253;
// bram[61607] = 251;
// bram[61608] = 244;
// bram[61609] = 232;
// bram[61610] = 215;
// bram[61611] = 195;
// bram[61612] = 172;
// bram[61613] = 146;
// bram[61614] = 120;
// bram[61615] = 95;
// bram[61616] = 70;
// bram[61617] = 48;
// bram[61618] = 29;
// bram[61619] = 15;
// bram[61620] = 5;
// bram[61621] = 0;
// bram[61622] = 0;
// bram[61623] = 6;
// bram[61624] = 17;
// bram[61625] = 32;
// bram[61626] = 52;
// bram[61627] = 74;
// bram[61628] = 99;
// bram[61629] = 125;
// bram[61630] = 151;
// bram[61631] = 176;
// bram[61632] = 199;
// bram[61633] = 218;
// bram[61634] = 234;
// bram[61635] = 246;
// bram[61636] = 252;
// bram[61637] = 253;
// bram[61638] = 249;
// bram[61639] = 240;
// bram[61640] = 226;
// bram[61641] = 207;
// bram[61642] = 186;
// bram[61643] = 162;
// bram[61644] = 136;
// bram[61645] = 110;
// bram[61646] = 85;
// bram[61647] = 61;
// bram[61648] = 40;
// bram[61649] = 23;
// bram[61650] = 10;
// bram[61651] = 2;
// bram[61652] = 0;
// bram[61653] = 2;
// bram[61654] = 10;
// bram[61655] = 23;
// bram[61656] = 40;
// bram[61657] = 61;
// bram[61658] = 84;
// bram[61659] = 109;
// bram[61660] = 135;
// bram[61661] = 161;
// bram[61662] = 185;
// bram[61663] = 207;
// bram[61664] = 225;
// bram[61665] = 240;
// bram[61666] = 249;
// bram[61667] = 253;
// bram[61668] = 252;
// bram[61669] = 246;
// bram[61670] = 235;
// bram[61671] = 219;
// bram[61672] = 199;
// bram[61673] = 176;
// bram[61674] = 151;
// bram[61675] = 125;
// bram[61676] = 99;
// bram[61677] = 75;
// bram[61678] = 52;
// bram[61679] = 33;
// bram[61680] = 17;
// bram[61681] = 6;
// bram[61682] = 0;
// bram[61683] = 0;
// bram[61684] = 5;
// bram[61685] = 15;
// bram[61686] = 29;
// bram[61687] = 48;
// bram[61688] = 70;
// bram[61689] = 94;
// bram[61690] = 120;
// bram[61691] = 146;
// bram[61692] = 171;
// bram[61693] = 195;
// bram[61694] = 215;
// bram[61695] = 232;
// bram[61696] = 244;
// bram[61697] = 251;
// bram[61698] = 253;
// bram[61699] = 250;
// bram[61700] = 242;
// bram[61701] = 229;
// bram[61702] = 211;
// bram[61703] = 190;
// bram[61704] = 166;
// bram[61705] = 141;
// bram[61706] = 115;
// bram[61707] = 89;
// bram[61708] = 65;
// bram[61709] = 44;
// bram[61710] = 26;
// bram[61711] = 12;
// bram[61712] = 3;
// bram[61713] = 0;
// bram[61714] = 1;
// bram[61715] = 8;
// bram[61716] = 20;
// bram[61717] = 36;
// bram[61718] = 57;
// bram[61719] = 80;
// bram[61720] = 105;
// bram[61721] = 131;
// bram[61722] = 156;
// bram[61723] = 181;
// bram[61724] = 203;
// bram[61725] = 222;
// bram[61726] = 237;
// bram[61727] = 248;
// bram[61728] = 253;
// bram[61729] = 253;
// bram[61730] = 247;
// bram[61731] = 237;
// bram[61732] = 222;
// bram[61733] = 203;
// bram[61734] = 180;
// bram[61735] = 156;
// bram[61736] = 130;
// bram[61737] = 104;
// bram[61738] = 79;
// bram[61739] = 56;
// bram[61740] = 36;
// bram[61741] = 20;
// bram[61742] = 8;
// bram[61743] = 1;
// bram[61744] = 0;
// bram[61745] = 3;
// bram[61746] = 12;
// bram[61747] = 26;
// bram[61748] = 44;
// bram[61749] = 66;
// bram[61750] = 90;
// bram[61751] = 115;
// bram[61752] = 141;
// bram[61753] = 167;
// bram[61754] = 190;
// bram[61755] = 211;
// bram[61756] = 229;
// bram[61757] = 242;
// bram[61758] = 250;
// bram[61759] = 253;
// bram[61760] = 251;
// bram[61761] = 244;
// bram[61762] = 231;
// bram[61763] = 215;
// bram[61764] = 194;
// bram[61765] = 171;
// bram[61766] = 145;
// bram[61767] = 119;
// bram[61768] = 94;
// bram[61769] = 69;
// bram[61770] = 47;
// bram[61771] = 29;
// bram[61772] = 14;
// bram[61773] = 5;
// bram[61774] = 0;
// bram[61775] = 1;
// bram[61776] = 6;
// bram[61777] = 17;
// bram[61778] = 33;
// bram[61779] = 53;
// bram[61780] = 75;
// bram[61781] = 100;
// bram[61782] = 126;
// bram[61783] = 152;
// bram[61784] = 177;
// bram[61785] = 199;
// bram[61786] = 219;
// bram[61787] = 235;
// bram[61788] = 246;
// bram[61789] = 252;
// bram[61790] = 253;
// bram[61791] = 249;
// bram[61792] = 239;
// bram[61793] = 225;
// bram[61794] = 207;
// bram[61795] = 185;
// bram[61796] = 161;
// bram[61797] = 135;
// bram[61798] = 109;
// bram[61799] = 84;
// bram[61800] = 60;
// bram[61801] = 39;
// bram[61802] = 22;
// bram[61803] = 10;
// bram[61804] = 2;
// bram[61805] = 0;
// bram[61806] = 2;
// bram[61807] = 10;
// bram[61808] = 23;
// bram[61809] = 41;
// bram[61810] = 61;
// bram[61811] = 85;
// bram[61812] = 110;
// bram[61813] = 136;
// bram[61814] = 162;
// bram[61815] = 186;
// bram[61816] = 208;
// bram[61817] = 226;
// bram[61818] = 240;
// bram[61819] = 249;
// bram[61820] = 253;
// bram[61821] = 252;
// bram[61822] = 246;
// bram[61823] = 234;
// bram[61824] = 218;
// bram[61825] = 198;
// bram[61826] = 175;
// bram[61827] = 150;
// bram[61828] = 124;
// bram[61829] = 98;
// bram[61830] = 74;
// bram[61831] = 51;
// bram[61832] = 32;
// bram[61833] = 17;
// bram[61834] = 6;
// bram[61835] = 0;
// bram[61836] = 0;
// bram[61837] = 5;
// bram[61838] = 15;
// bram[61839] = 30;
// bram[61840] = 49;
// bram[61841] = 71;
// bram[61842] = 95;
// bram[61843] = 121;
// bram[61844] = 147;
// bram[61845] = 172;
// bram[61846] = 195;
// bram[61847] = 216;
// bram[61848] = 232;
// bram[61849] = 244;
// bram[61850] = 252;
// bram[61851] = 253;
// bram[61852] = 250;
// bram[61853] = 241;
// bram[61854] = 228;
// bram[61855] = 210;
// bram[61856] = 189;
// bram[61857] = 165;
// bram[61858] = 140;
// bram[61859] = 114;
// bram[61860] = 88;
// bram[61861] = 64;
// bram[61862] = 43;
// bram[61863] = 25;
// bram[61864] = 12;
// bram[61865] = 3;
// bram[61866] = 0;
// bram[61867] = 1;
// bram[61868] = 8;
// bram[61869] = 21;
// bram[61870] = 37;
// bram[61871] = 57;
// bram[61872] = 80;
// bram[61873] = 106;
// bram[61874] = 132;
// bram[61875] = 157;
// bram[61876] = 182;
// bram[61877] = 204;
// bram[61878] = 223;
// bram[61879] = 238;
// bram[61880] = 248;
// bram[61881] = 253;
// bram[61882] = 253;
// bram[61883] = 247;
// bram[61884] = 237;
// bram[61885] = 221;
// bram[61886] = 202;
// bram[61887] = 180;
// bram[61888] = 155;
// bram[61889] = 129;
// bram[61890] = 103;
// bram[61891] = 78;
// bram[61892] = 55;
// bram[61893] = 35;
// bram[61894] = 19;
// bram[61895] = 8;
// bram[61896] = 1;
// bram[61897] = 0;
// bram[61898] = 4;
// bram[61899] = 13;
// bram[61900] = 27;
// bram[61901] = 45;
// bram[61902] = 66;
// bram[61903] = 91;
// bram[61904] = 116;
// bram[61905] = 142;
// bram[61906] = 168;
// bram[61907] = 191;
// bram[61908] = 212;
// bram[61909] = 229;
// bram[61910] = 242;
// bram[61911] = 251;
// bram[61912] = 253;
// bram[61913] = 251;
// bram[61914] = 243;
// bram[61915] = 231;
// bram[61916] = 214;
// bram[61917] = 193;
// bram[61918] = 170;
// bram[61919] = 145;
// bram[61920] = 119;
// bram[61921] = 93;
// bram[61922] = 69;
// bram[61923] = 47;
// bram[61924] = 28;
// bram[61925] = 14;
// bram[61926] = 4;
// bram[61927] = 0;
// bram[61928] = 1;
// bram[61929] = 7;
// bram[61930] = 18;
// bram[61931] = 34;
// bram[61932] = 53;
// bram[61933] = 76;
// bram[61934] = 101;
// bram[61935] = 127;
// bram[61936] = 153;
// bram[61937] = 177;
// bram[61938] = 200;
// bram[61939] = 220;
// bram[61940] = 235;
// bram[61941] = 246;
// bram[61942] = 252;
// bram[61943] = 253;
// bram[61944] = 249;
// bram[61945] = 239;
// bram[61946] = 224;
// bram[61947] = 206;
// bram[61948] = 184;
// bram[61949] = 160;
// bram[61950] = 134;
// bram[61951] = 108;
// bram[61952] = 83;
// bram[61953] = 59;
// bram[61954] = 39;
// bram[61955] = 22;
// bram[61956] = 9;
// bram[61957] = 2;
// bram[61958] = 0;
// bram[61959] = 3;
// bram[61960] = 11;
// bram[61961] = 24;
// bram[61962] = 41;
// bram[61963] = 62;
// bram[61964] = 86;
// bram[61965] = 111;
// bram[61966] = 137;
// bram[61967] = 163;
// bram[61968] = 187;
// bram[61969] = 208;
// bram[61970] = 227;
// bram[61971] = 240;
// bram[61972] = 249;
// bram[61973] = 253;
// bram[61974] = 252;
// bram[61975] = 245;
// bram[61976] = 234;
// bram[61977] = 217;
// bram[61978] = 197;
// bram[61979] = 174;
// bram[61980] = 149;
// bram[61981] = 123;
// bram[61982] = 98;
// bram[61983] = 73;
// bram[61984] = 51;
// bram[61985] = 31;
// bram[61986] = 16;
// bram[61987] = 6;
// bram[61988] = 0;
// bram[61989] = 0;
// bram[61990] = 5;
// bram[61991] = 16;
// bram[61992] = 30;
// bram[61993] = 49;
// bram[61994] = 72;
// bram[61995] = 96;
// bram[61996] = 122;
// bram[61997] = 148;
// bram[61998] = 173;
// bram[61999] = 196;
// bram[62000] = 216;
// bram[62001] = 233;
// bram[62002] = 245;
// bram[62003] = 252;
// bram[62004] = 253;
// bram[62005] = 250;
// bram[62006] = 241;
// bram[62007] = 227;
// bram[62008] = 210;
// bram[62009] = 188;
// bram[62010] = 164;
// bram[62011] = 139;
// bram[62012] = 113;
// bram[62013] = 87;
// bram[62014] = 63;
// bram[62015] = 42;
// bram[62016] = 25;
// bram[62017] = 11;
// bram[62018] = 3;
// bram[62019] = 0;
// bram[62020] = 2;
// bram[62021] = 9;
// bram[62022] = 21;
// bram[62023] = 38;
// bram[62024] = 58;
// bram[62025] = 81;
// bram[62026] = 107;
// bram[62027] = 133;
// bram[62028] = 158;
// bram[62029] = 183;
// bram[62030] = 205;
// bram[62031] = 223;
// bram[62032] = 238;
// bram[62033] = 248;
// bram[62034] = 253;
// bram[62035] = 253;
// bram[62036] = 247;
// bram[62037] = 236;
// bram[62038] = 221;
// bram[62039] = 201;
// bram[62040] = 179;
// bram[62041] = 154;
// bram[62042] = 128;
// bram[62043] = 102;
// bram[62044] = 77;
// bram[62045] = 54;
// bram[62046] = 35;
// bram[62047] = 19;
// bram[62048] = 7;
// bram[62049] = 1;
// bram[62050] = 0;
// bram[62051] = 4;
// bram[62052] = 13;
// bram[62053] = 27;
// bram[62054] = 46;
// bram[62055] = 67;
// bram[62056] = 91;
// bram[62057] = 117;
// bram[62058] = 143;
// bram[62059] = 168;
// bram[62060] = 192;
// bram[62061] = 213;
// bram[62062] = 230;
// bram[62063] = 243;
// bram[62064] = 251;
// bram[62065] = 253;
// bram[62066] = 251;
// bram[62067] = 243;
// bram[62068] = 230;
// bram[62069] = 213;
// bram[62070] = 192;
// bram[62071] = 169;
// bram[62072] = 144;
// bram[62073] = 118;
// bram[62074] = 92;
// bram[62075] = 68;
// bram[62076] = 46;
// bram[62077] = 28;
// bram[62078] = 13;
// bram[62079] = 4;
// bram[62080] = 0;
// bram[62081] = 1;
// bram[62082] = 7;
// bram[62083] = 18;
// bram[62084] = 34;
// bram[62085] = 54;
// bram[62086] = 77;
// bram[62087] = 102;
// bram[62088] = 128;
// bram[62089] = 154;
// bram[62090] = 178;
// bram[62091] = 201;
// bram[62092] = 220;
// bram[62093] = 236;
// bram[62094] = 247;
// bram[62095] = 253;
// bram[62096] = 253;
// bram[62097] = 248;
// bram[62098] = 238;
// bram[62099] = 224;
// bram[62100] = 205;
// bram[62101] = 183;
// bram[62102] = 159;
// bram[62103] = 133;
// bram[62104] = 107;
// bram[62105] = 82;
// bram[62106] = 59;
// bram[62107] = 38;
// bram[62108] = 21;
// bram[62109] = 9;
// bram[62110] = 2;
// bram[62111] = 0;
// bram[62112] = 3;
// bram[62113] = 11;
// bram[62114] = 24;
// bram[62115] = 42;
// bram[62116] = 63;
// bram[62117] = 87;
// bram[62118] = 112;
// bram[62119] = 138;
// bram[62120] = 164;
// bram[62121] = 188;
// bram[62122] = 209;
// bram[62123] = 227;
// bram[62124] = 241;
// bram[62125] = 250;
// bram[62126] = 253;
// bram[62127] = 252;
// bram[62128] = 245;
// bram[62129] = 233;
// bram[62130] = 217;
// bram[62131] = 197;
// bram[62132] = 173;
// bram[62133] = 148;
// bram[62134] = 122;
// bram[62135] = 97;
// bram[62136] = 72;
// bram[62137] = 50;
// bram[62138] = 31;
// bram[62139] = 16;
// bram[62140] = 5;
// bram[62141] = 0;
// bram[62142] = 0;
// bram[62143] = 6;
// bram[62144] = 16;
// bram[62145] = 31;
// bram[62146] = 50;
// bram[62147] = 72;
// bram[62148] = 97;
// bram[62149] = 123;
// bram[62150] = 149;
// bram[62151] = 174;
// bram[62152] = 197;
// bram[62153] = 217;
// bram[62154] = 233;
// bram[62155] = 245;
// bram[62156] = 252;
// bram[62157] = 253;
// bram[62158] = 250;
// bram[62159] = 241;
// bram[62160] = 227;
// bram[62161] = 209;
// bram[62162] = 187;
// bram[62163] = 163;
// bram[62164] = 138;
// bram[62165] = 112;
// bram[62166] = 86;
// bram[62167] = 63;
// bram[62168] = 42;
// bram[62169] = 24;
// bram[62170] = 11;
// bram[62171] = 3;
// bram[62172] = 0;
// bram[62173] = 2;
// bram[62174] = 9;
// bram[62175] = 22;
// bram[62176] = 38;
// bram[62177] = 59;
// bram[62178] = 82;
// bram[62179] = 107;
// bram[62180] = 133;
// bram[62181] = 159;
// bram[62182] = 184;
// bram[62183] = 205;
// bram[62184] = 224;
// bram[62185] = 239;
// bram[62186] = 248;
// bram[62187] = 253;
// bram[62188] = 252;
// bram[62189] = 247;
// bram[62190] = 236;
// bram[62191] = 220;
// bram[62192] = 201;
// bram[62193] = 178;
// bram[62194] = 153;
// bram[62195] = 127;
// bram[62196] = 101;
// bram[62197] = 76;
// bram[62198] = 54;
// bram[62199] = 34;
// bram[62200] = 18;
// bram[62201] = 7;
// bram[62202] = 1;
// bram[62203] = 0;
// bram[62204] = 4;
// bram[62205] = 14;
// bram[62206] = 28;
// bram[62207] = 46;
// bram[62208] = 68;
// bram[62209] = 92;
// bram[62210] = 118;
// bram[62211] = 144;
// bram[62212] = 169;
// bram[62213] = 193;
// bram[62214] = 214;
// bram[62215] = 231;
// bram[62216] = 243;
// bram[62217] = 251;
// bram[62218] = 253;
// bram[62219] = 251;
// bram[62220] = 243;
// bram[62221] = 230;
// bram[62222] = 212;
// bram[62223] = 192;
// bram[62224] = 168;
// bram[62225] = 143;
// bram[62226] = 117;
// bram[62227] = 91;
// bram[62228] = 67;
// bram[62229] = 45;
// bram[62230] = 27;
// bram[62231] = 13;
// bram[62232] = 4;
// bram[62233] = 0;
// bram[62234] = 1;
// bram[62235] = 7;
// bram[62236] = 19;
// bram[62237] = 35;
// bram[62238] = 55;
// bram[62239] = 78;
// bram[62240] = 103;
// bram[62241] = 129;
// bram[62242] = 154;
// bram[62243] = 179;
// bram[62244] = 202;
// bram[62245] = 221;
// bram[62246] = 236;
// bram[62247] = 247;
// bram[62248] = 253;
// bram[62249] = 253;
// bram[62250] = 248;
// bram[62251] = 238;
// bram[62252] = 223;
// bram[62253] = 204;
// bram[62254] = 182;
// bram[62255] = 158;
// bram[62256] = 132;
// bram[62257] = 106;
// bram[62258] = 81;
// bram[62259] = 58;
// bram[62260] = 37;
// bram[62261] = 21;
// bram[62262] = 9;
// bram[62263] = 1;
// bram[62264] = 0;
// bram[62265] = 3;
// bram[62266] = 12;
// bram[62267] = 25;
// bram[62268] = 43;
// bram[62269] = 64;
// bram[62270] = 88;
// bram[62271] = 113;
// bram[62272] = 139;
// bram[62273] = 165;
// bram[62274] = 189;
// bram[62275] = 210;
// bram[62276] = 228;
// bram[62277] = 241;
// bram[62278] = 250;
// bram[62279] = 253;
// bram[62280] = 252;
// bram[62281] = 245;
// bram[62282] = 232;
// bram[62283] = 216;
// bram[62284] = 196;
// bram[62285] = 173;
// bram[62286] = 147;
// bram[62287] = 121;
// bram[62288] = 96;
// bram[62289] = 71;
// bram[62290] = 49;
// bram[62291] = 30;
// bram[62292] = 15;
// bram[62293] = 5;
// bram[62294] = 0;
// bram[62295] = 0;
// bram[62296] = 6;
// bram[62297] = 16;
// bram[62298] = 32;
// bram[62299] = 51;
// bram[62300] = 73;
// bram[62301] = 98;
// bram[62302] = 124;
// bram[62303] = 150;
// bram[62304] = 175;
// bram[62305] = 198;
// bram[62306] = 218;
// bram[62307] = 234;
// bram[62308] = 245;
// bram[62309] = 252;
// bram[62310] = 253;
// bram[62311] = 249;
// bram[62312] = 240;
// bram[62313] = 226;
// bram[62314] = 208;
// bram[62315] = 187;
// bram[62316] = 163;
// bram[62317] = 137;
// bram[62318] = 111;
// bram[62319] = 86;
// bram[62320] = 62;
// bram[62321] = 41;
// bram[62322] = 24;
// bram[62323] = 11;
// bram[62324] = 2;
// bram[62325] = 0;
// bram[62326] = 2;
// bram[62327] = 10;
// bram[62328] = 22;
// bram[62329] = 39;
// bram[62330] = 60;
// bram[62331] = 83;
// bram[62332] = 108;
// bram[62333] = 134;
// bram[62334] = 160;
// bram[62335] = 184;
// bram[62336] = 206;
// bram[62337] = 225;
// bram[62338] = 239;
// bram[62339] = 249;
// bram[62340] = 253;
// bram[62341] = 252;
// bram[62342] = 246;
// bram[62343] = 235;
// bram[62344] = 219;
// bram[62345] = 200;
// bram[62346] = 177;
// bram[62347] = 152;
// bram[62348] = 126;
// bram[62349] = 100;
// bram[62350] = 76;
// bram[62351] = 53;
// bram[62352] = 33;
// bram[62353] = 18;
// bram[62354] = 7;
// bram[62355] = 1;
// bram[62356] = 0;
// bram[62357] = 4;
// bram[62358] = 14;
// bram[62359] = 29;
// bram[62360] = 47;
// bram[62361] = 69;
// bram[62362] = 93;
// bram[62363] = 119;
// bram[62364] = 145;
// bram[62365] = 170;
// bram[62366] = 194;
// bram[62367] = 214;
// bram[62368] = 231;
// bram[62369] = 244;
// bram[62370] = 251;
// bram[62371] = 253;
// bram[62372] = 250;
// bram[62373] = 242;
// bram[62374] = 229;
// bram[62375] = 212;
// bram[62376] = 191;
// bram[62377] = 167;
// bram[62378] = 142;
// bram[62379] = 116;
// bram[62380] = 90;
// bram[62381] = 66;
// bram[62382] = 45;
// bram[62383] = 26;
// bram[62384] = 13;
// bram[62385] = 4;
// bram[62386] = 0;
// bram[62387] = 1;
// bram[62388] = 8;
// bram[62389] = 19;
// bram[62390] = 36;
// bram[62391] = 56;
// bram[62392] = 79;
// bram[62393] = 104;
// bram[62394] = 130;
// bram[62395] = 155;
// bram[62396] = 180;
// bram[62397] = 202;
// bram[62398] = 222;
// bram[62399] = 237;
// bram[62400] = 247;
// bram[62401] = 253;
// bram[62402] = 253;
// bram[62403] = 248;
// bram[62404] = 238;
// bram[62405] = 223;
// bram[62406] = 204;
// bram[62407] = 181;
// bram[62408] = 157;
// bram[62409] = 131;
// bram[62410] = 105;
// bram[62411] = 80;
// bram[62412] = 57;
// bram[62413] = 37;
// bram[62414] = 20;
// bram[62415] = 8;
// bram[62416] = 1;
// bram[62417] = 0;
// bram[62418] = 3;
// bram[62419] = 12;
// bram[62420] = 26;
// bram[62421] = 43;
// bram[62422] = 65;
// bram[62423] = 89;
// bram[62424] = 114;
// bram[62425] = 140;
// bram[62426] = 166;
// bram[62427] = 189;
// bram[62428] = 211;
// bram[62429] = 228;
// bram[62430] = 242;
// bram[62431] = 250;
// bram[62432] = 253;
// bram[62433] = 251;
// bram[62434] = 244;
// bram[62435] = 232;
// bram[62436] = 215;
// bram[62437] = 195;
// bram[62438] = 172;
// bram[62439] = 147;
// bram[62440] = 121;
// bram[62441] = 95;
// bram[62442] = 70;
// bram[62443] = 48;
// bram[62444] = 30;
// bram[62445] = 15;
// bram[62446] = 5;
// bram[62447] = 0;
// bram[62448] = 0;
// bram[62449] = 6;
// bram[62450] = 17;
// bram[62451] = 32;
// bram[62452] = 52;
// bram[62453] = 74;
// bram[62454] = 99;
// bram[62455] = 125;
// bram[62456] = 151;
// bram[62457] = 176;
// bram[62458] = 198;
// bram[62459] = 218;
// bram[62460] = 234;
// bram[62461] = 246;
// bram[62462] = 252;
// bram[62463] = 253;
// bram[62464] = 249;
// bram[62465] = 240;
// bram[62466] = 226;
// bram[62467] = 207;
// bram[62468] = 186;
// bram[62469] = 162;
// bram[62470] = 136;
// bram[62471] = 110;
// bram[62472] = 85;
// bram[62473] = 61;
// bram[62474] = 40;
// bram[62475] = 23;
// bram[62476] = 10;
// bram[62477] = 2;
// bram[62478] = 0;
// bram[62479] = 2;
// bram[62480] = 10;
// bram[62481] = 23;
// bram[62482] = 40;
// bram[62483] = 61;
// bram[62484] = 84;
// bram[62485] = 109;
// bram[62486] = 135;
// bram[62487] = 161;
// bram[62488] = 185;
// bram[62489] = 207;
// bram[62490] = 225;
// bram[62491] = 239;
// bram[62492] = 249;
// bram[62493] = 253;
// bram[62494] = 252;
// bram[62495] = 246;
// bram[62496] = 235;
// bram[62497] = 219;
// bram[62498] = 199;
// bram[62499] = 176;
// bram[62500] = 151;
// bram[62501] = 125;
// bram[62502] = 99;
// bram[62503] = 75;
// bram[62504] = 52;
// bram[62505] = 33;
// bram[62506] = 17;
// bram[62507] = 6;
// bram[62508] = 0;
// bram[62509] = 0;
// bram[62510] = 5;
// bram[62511] = 15;
// bram[62512] = 29;
// bram[62513] = 48;
// bram[62514] = 70;
// bram[62515] = 94;
// bram[62516] = 120;
// bram[62517] = 146;
// bram[62518] = 171;
// bram[62519] = 194;
// bram[62520] = 215;
// bram[62521] = 232;
// bram[62522] = 244;
// bram[62523] = 251;
// bram[62524] = 253;
// bram[62525] = 250;
// bram[62526] = 242;
// bram[62527] = 229;
// bram[62528] = 211;
// bram[62529] = 190;
// bram[62530] = 166;
// bram[62531] = 141;
// bram[62532] = 115;
// bram[62533] = 89;
// bram[62534] = 65;
// bram[62535] = 44;
// bram[62536] = 26;
// bram[62537] = 12;
// bram[62538] = 3;
// bram[62539] = 0;
// bram[62540] = 1;
// bram[62541] = 8;
// bram[62542] = 20;
// bram[62543] = 36;
// bram[62544] = 56;
// bram[62545] = 80;
// bram[62546] = 105;
// bram[62547] = 131;
// bram[62548] = 156;
// bram[62549] = 181;
// bram[62550] = 203;
// bram[62551] = 222;
// bram[62552] = 237;
// bram[62553] = 248;
// bram[62554] = 253;
// bram[62555] = 253;
// bram[62556] = 247;
// bram[62557] = 237;
// bram[62558] = 222;
// bram[62559] = 203;
// bram[62560] = 181;
// bram[62561] = 156;
// bram[62562] = 130;
// bram[62563] = 104;
// bram[62564] = 79;
// bram[62565] = 56;
// bram[62566] = 36;
// bram[62567] = 20;
// bram[62568] = 8;
// bram[62569] = 1;
// bram[62570] = 0;
// bram[62571] = 3;
// bram[62572] = 12;
// bram[62573] = 26;
// bram[62574] = 44;
// bram[62575] = 66;
// bram[62576] = 90;
// bram[62577] = 115;
// bram[62578] = 141;
// bram[62579] = 167;
// bram[62580] = 190;
// bram[62581] = 211;
// bram[62582] = 229;
// bram[62583] = 242;
// bram[62584] = 250;
// bram[62585] = 253;
// bram[62586] = 251;
// bram[62587] = 244;
// bram[62588] = 231;
// bram[62589] = 215;
// bram[62590] = 194;
// bram[62591] = 171;
// bram[62592] = 146;
// bram[62593] = 120;
// bram[62594] = 94;
// bram[62595] = 70;
// bram[62596] = 48;
// bram[62597] = 29;
// bram[62598] = 14;
// bram[62599] = 5;
// bram[62600] = 0;
// bram[62601] = 1;
// bram[62602] = 6;
// bram[62603] = 17;
// bram[62604] = 33;
// bram[62605] = 52;
// bram[62606] = 75;
// bram[62607] = 100;
// bram[62608] = 126;
// bram[62609] = 152;
// bram[62610] = 176;
// bram[62611] = 199;
// bram[62612] = 219;
// bram[62613] = 235;
// bram[62614] = 246;
// bram[62615] = 252;
// bram[62616] = 253;
// bram[62617] = 249;
// bram[62618] = 239;
// bram[62619] = 225;
// bram[62620] = 207;
// bram[62621] = 185;
// bram[62622] = 161;
// bram[62623] = 135;
// bram[62624] = 109;
// bram[62625] = 84;
// bram[62626] = 60;
// bram[62627] = 40;
// bram[62628] = 22;
// bram[62629] = 10;
// bram[62630] = 2;
// bram[62631] = 0;
// bram[62632] = 2;
// bram[62633] = 10;
// bram[62634] = 23;
// bram[62635] = 40;
// bram[62636] = 61;
// bram[62637] = 85;
// bram[62638] = 110;
// bram[62639] = 136;
// bram[62640] = 162;
// bram[62641] = 186;
// bram[62642] = 208;
// bram[62643] = 226;
// bram[62644] = 240;
// bram[62645] = 249;
// bram[62646] = 253;
// bram[62647] = 252;
// bram[62648] = 246;
// bram[62649] = 234;
// bram[62650] = 218;
// bram[62651] = 198;
// bram[62652] = 175;
// bram[62653] = 150;
// bram[62654] = 124;
// bram[62655] = 99;
// bram[62656] = 74;
// bram[62657] = 51;
// bram[62658] = 32;
// bram[62659] = 17;
// bram[62660] = 6;
// bram[62661] = 0;
// bram[62662] = 0;
// bram[62663] = 5;
// bram[62664] = 15;
// bram[62665] = 30;
// bram[62666] = 49;
// bram[62667] = 71;
// bram[62668] = 95;
// bram[62669] = 121;
// bram[62670] = 147;
// bram[62671] = 172;
// bram[62672] = 195;
// bram[62673] = 216;
// bram[62674] = 232;
// bram[62675] = 244;
// bram[62676] = 252;
// bram[62677] = 253;
// bram[62678] = 250;
// bram[62679] = 241;
// bram[62680] = 228;
// bram[62681] = 210;
// bram[62682] = 189;
// bram[62683] = 165;
// bram[62684] = 140;
// bram[62685] = 114;
// bram[62686] = 88;
// bram[62687] = 64;
// bram[62688] = 43;
// bram[62689] = 25;
// bram[62690] = 12;
// bram[62691] = 3;
// bram[62692] = 0;
// bram[62693] = 1;
// bram[62694] = 8;
// bram[62695] = 20;
// bram[62696] = 37;
// bram[62697] = 57;
// bram[62698] = 80;
// bram[62699] = 106;
// bram[62700] = 131;
// bram[62701] = 157;
// bram[62702] = 182;
// bram[62703] = 204;
// bram[62704] = 223;
// bram[62705] = 238;
// bram[62706] = 248;
// bram[62707] = 253;
// bram[62708] = 253;
// bram[62709] = 247;
// bram[62710] = 237;
// bram[62711] = 221;
// bram[62712] = 202;
// bram[62713] = 180;
// bram[62714] = 155;
// bram[62715] = 129;
// bram[62716] = 103;
// bram[62717] = 78;
// bram[62718] = 55;
// bram[62719] = 35;
// bram[62720] = 19;
// bram[62721] = 8;
// bram[62722] = 1;
// bram[62723] = 0;
// bram[62724] = 4;
// bram[62725] = 13;
// bram[62726] = 27;
// bram[62727] = 45;
// bram[62728] = 66;
// bram[62729] = 90;
// bram[62730] = 116;
// bram[62731] = 142;
// bram[62732] = 167;
// bram[62733] = 191;
// bram[62734] = 212;
// bram[62735] = 229;
// bram[62736] = 242;
// bram[62737] = 251;
// bram[62738] = 253;
// bram[62739] = 251;
// bram[62740] = 243;
// bram[62741] = 231;
// bram[62742] = 214;
// bram[62743] = 193;
// bram[62744] = 170;
// bram[62745] = 145;
// bram[62746] = 119;
// bram[62747] = 93;
// bram[62748] = 69;
// bram[62749] = 47;
// bram[62750] = 28;
// bram[62751] = 14;
// bram[62752] = 4;
// bram[62753] = 0;
// bram[62754] = 1;
// bram[62755] = 7;
// bram[62756] = 18;
// bram[62757] = 34;
// bram[62758] = 53;
// bram[62759] = 76;
// bram[62760] = 101;
// bram[62761] = 127;
// bram[62762] = 153;
// bram[62763] = 177;
// bram[62764] = 200;
// bram[62765] = 220;
// bram[62766] = 235;
// bram[62767] = 246;
// bram[62768] = 252;
// bram[62769] = 253;
// bram[62770] = 249;
// bram[62771] = 239;
// bram[62772] = 224;
// bram[62773] = 206;
// bram[62774] = 184;
// bram[62775] = 160;
// bram[62776] = 134;
// bram[62777] = 108;
// bram[62778] = 83;
// bram[62779] = 59;
// bram[62780] = 39;
// bram[62781] = 22;
// bram[62782] = 9;
// bram[62783] = 2;
// bram[62784] = 0;
// bram[62785] = 3;
// bram[62786] = 11;
// bram[62787] = 24;
// bram[62788] = 41;
// bram[62789] = 62;
// bram[62790] = 86;
// bram[62791] = 111;
// bram[62792] = 137;
// bram[62793] = 163;
// bram[62794] = 187;
// bram[62795] = 208;
// bram[62796] = 226;
// bram[62797] = 240;
// bram[62798] = 249;
// bram[62799] = 253;
// bram[62800] = 252;
// bram[62801] = 245;
// bram[62802] = 234;
// bram[62803] = 217;
// bram[62804] = 197;
// bram[62805] = 174;
// bram[62806] = 149;
// bram[62807] = 123;
// bram[62808] = 98;
// bram[62809] = 73;
// bram[62810] = 51;
// bram[62811] = 31;
// bram[62812] = 16;
// bram[62813] = 6;
// bram[62814] = 0;
// bram[62815] = 0;
// bram[62816] = 5;
// bram[62817] = 15;
// bram[62818] = 30;
// bram[62819] = 49;
// bram[62820] = 72;
// bram[62821] = 96;
// bram[62822] = 122;
// bram[62823] = 148;
// bram[62824] = 173;
// bram[62825] = 196;
// bram[62826] = 216;
// bram[62827] = 233;
// bram[62828] = 245;
// bram[62829] = 252;
// bram[62830] = 253;
// bram[62831] = 250;
// bram[62832] = 241;
// bram[62833] = 227;
// bram[62834] = 210;
// bram[62835] = 188;
// bram[62836] = 164;
// bram[62837] = 139;
// bram[62838] = 113;
// bram[62839] = 87;
// bram[62840] = 64;
// bram[62841] = 42;
// bram[62842] = 25;
// bram[62843] = 11;
// bram[62844] = 3;
// bram[62845] = 0;
// bram[62846] = 2;
// bram[62847] = 9;
// bram[62848] = 21;
// bram[62849] = 38;
// bram[62850] = 58;
// bram[62851] = 81;
// bram[62852] = 106;
// bram[62853] = 132;
// bram[62854] = 158;
// bram[62855] = 183;
// bram[62856] = 205;
// bram[62857] = 223;
// bram[62858] = 238;
// bram[62859] = 248;
// bram[62860] = 253;
// bram[62861] = 253;
// bram[62862] = 247;
// bram[62863] = 236;
// bram[62864] = 221;
// bram[62865] = 201;
// bram[62866] = 179;
// bram[62867] = 154;
// bram[62868] = 128;
// bram[62869] = 102;
// bram[62870] = 77;
// bram[62871] = 55;
// bram[62872] = 35;
// bram[62873] = 19;
// bram[62874] = 7;
// bram[62875] = 1;
// bram[62876] = 0;
// bram[62877] = 4;
// bram[62878] = 13;
// bram[62879] = 27;
// bram[62880] = 46;
// bram[62881] = 67;
// bram[62882] = 91;
// bram[62883] = 117;
// bram[62884] = 143;
// bram[62885] = 168;
// bram[62886] = 192;
// bram[62887] = 213;
// bram[62888] = 230;
// bram[62889] = 243;
// bram[62890] = 251;
// bram[62891] = 253;
// bram[62892] = 251;
// bram[62893] = 243;
// bram[62894] = 230;
// bram[62895] = 213;
// bram[62896] = 193;
// bram[62897] = 169;
// bram[62898] = 144;
// bram[62899] = 118;
// bram[62900] = 92;
// bram[62901] = 68;
// bram[62902] = 46;
// bram[62903] = 28;
// bram[62904] = 14;
// bram[62905] = 4;
// bram[62906] = 0;
// bram[62907] = 1;
// bram[62908] = 7;
// bram[62909] = 18;
// bram[62910] = 34;
// bram[62911] = 54;
// bram[62912] = 77;
// bram[62913] = 102;
// bram[62914] = 128;
// bram[62915] = 153;
// bram[62916] = 178;
// bram[62917] = 201;
// bram[62918] = 220;
// bram[62919] = 236;
// bram[62920] = 247;
// bram[62921] = 253;
// bram[62922] = 253;
// bram[62923] = 248;
// bram[62924] = 238;
// bram[62925] = 224;
// bram[62926] = 205;
// bram[62927] = 183;
// bram[62928] = 159;
// bram[62929] = 133;
// bram[62930] = 107;
// bram[62931] = 82;
// bram[62932] = 59;
// bram[62933] = 38;
// bram[62934] = 21;
// bram[62935] = 9;
// bram[62936] = 2;
// bram[62937] = 0;
// bram[62938] = 3;
// bram[62939] = 11;
// bram[62940] = 24;
// bram[62941] = 42;
// bram[62942] = 63;
// bram[62943] = 87;
// bram[62944] = 112;
// bram[62945] = 138;
// bram[62946] = 164;
// bram[62947] = 188;
// bram[62948] = 209;
// bram[62949] = 227;
// bram[62950] = 241;
// bram[62951] = 250;
// bram[62952] = 253;
// bram[62953] = 252;
// bram[62954] = 245;
// bram[62955] = 233;
// bram[62956] = 217;
// bram[62957] = 197;
// bram[62958] = 174;
// bram[62959] = 148;
// bram[62960] = 123;
// bram[62961] = 97;
// bram[62962] = 72;
// bram[62963] = 50;
// bram[62964] = 31;
// bram[62965] = 16;
// bram[62966] = 5;
// bram[62967] = 0;
// bram[62968] = 0;
// bram[62969] = 6;
// bram[62970] = 16;
// bram[62971] = 31;
// bram[62972] = 50;
// bram[62973] = 72;
// bram[62974] = 97;
// bram[62975] = 123;
// bram[62976] = 149;
// bram[62977] = 174;
// bram[62978] = 197;
// bram[62979] = 217;
// bram[62980] = 233;
// bram[62981] = 245;
// bram[62982] = 252;
// bram[62983] = 253;
// bram[62984] = 250;
// bram[62985] = 241;
// bram[62986] = 227;
// bram[62987] = 209;
// bram[62988] = 188;
// bram[62989] = 164;
// bram[62990] = 138;
// bram[62991] = 112;
// bram[62992] = 86;
// bram[62993] = 63;
// bram[62994] = 42;
// bram[62995] = 24;
// bram[62996] = 11;
// bram[62997] = 3;
// bram[62998] = 0;
// bram[62999] = 2;
// bram[63000] = 9;
// bram[63001] = 22;
// bram[63002] = 38;
// bram[63003] = 59;
// bram[63004] = 82;
// bram[63005] = 107;
// bram[63006] = 133;
// bram[63007] = 159;
// bram[63008] = 183;
// bram[63009] = 205;
// bram[63010] = 224;
// bram[63011] = 239;
// bram[63012] = 248;
// bram[63013] = 253;
// bram[63014] = 252;
// bram[63015] = 247;
// bram[63016] = 236;
// bram[63017] = 220;
// bram[63018] = 201;
// bram[63019] = 178;
// bram[63020] = 153;
// bram[63021] = 127;
// bram[63022] = 101;
// bram[63023] = 77;
// bram[63024] = 54;
// bram[63025] = 34;
// bram[63026] = 18;
// bram[63027] = 7;
// bram[63028] = 1;
// bram[63029] = 0;
// bram[63030] = 4;
// bram[63031] = 14;
// bram[63032] = 28;
// bram[63033] = 46;
// bram[63034] = 68;
// bram[63035] = 92;
// bram[63036] = 118;
// bram[63037] = 144;
// bram[63038] = 169;
// bram[63039] = 193;
// bram[63040] = 213;
// bram[63041] = 230;
// bram[63042] = 243;
// bram[63043] = 251;
// bram[63044] = 253;
// bram[63045] = 251;
// bram[63046] = 243;
// bram[63047] = 230;
// bram[63048] = 213;
// bram[63049] = 192;
// bram[63050] = 168;
// bram[63051] = 143;
// bram[63052] = 117;
// bram[63053] = 91;
// bram[63054] = 67;
// bram[63055] = 45;
// bram[63056] = 27;
// bram[63057] = 13;
// bram[63058] = 4;
// bram[63059] = 0;
// bram[63060] = 1;
// bram[63061] = 7;
// bram[63062] = 19;
// bram[63063] = 35;
// bram[63064] = 55;
// bram[63065] = 78;
// bram[63066] = 103;
// bram[63067] = 129;
// bram[63068] = 154;
// bram[63069] = 179;
// bram[63070] = 202;
// bram[63071] = 221;
// bram[63072] = 236;
// bram[63073] = 247;
// bram[63074] = 253;
// bram[63075] = 253;
// bram[63076] = 248;
// bram[63077] = 238;
// bram[63078] = 223;
// bram[63079] = 204;
// bram[63080] = 182;
// bram[63081] = 158;
// bram[63082] = 132;
// bram[63083] = 106;
// bram[63084] = 81;
// bram[63085] = 58;
// bram[63086] = 37;
// bram[63087] = 21;
// bram[63088] = 9;
// bram[63089] = 2;
// bram[63090] = 0;
// bram[63091] = 3;
// bram[63092] = 12;
// bram[63093] = 25;
// bram[63094] = 43;
// bram[63095] = 64;
// bram[63096] = 88;
// bram[63097] = 113;
// bram[63098] = 139;
// bram[63099] = 165;
// bram[63100] = 189;
// bram[63101] = 210;
// bram[63102] = 228;
// bram[63103] = 241;
// bram[63104] = 250;
// bram[63105] = 253;
// bram[63106] = 252;
// bram[63107] = 245;
// bram[63108] = 233;
// bram[63109] = 216;
// bram[63110] = 196;
// bram[63111] = 173;
// bram[63112] = 148;
// bram[63113] = 122;
// bram[63114] = 96;
// bram[63115] = 71;
// bram[63116] = 49;
// bram[63117] = 30;
// bram[63118] = 15;
// bram[63119] = 5;
// bram[63120] = 0;
// bram[63121] = 0;
// bram[63122] = 6;
// bram[63123] = 16;
// bram[63124] = 32;
// bram[63125] = 51;
// bram[63126] = 73;
// bram[63127] = 98;
// bram[63128] = 124;
// bram[63129] = 150;
// bram[63130] = 175;
// bram[63131] = 198;
// bram[63132] = 218;
// bram[63133] = 234;
// bram[63134] = 245;
// bram[63135] = 252;
// bram[63136] = 253;
// bram[63137] = 249;
// bram[63138] = 240;
// bram[63139] = 226;
// bram[63140] = 208;
// bram[63141] = 187;
// bram[63142] = 163;
// bram[63143] = 137;
// bram[63144] = 111;
// bram[63145] = 86;
// bram[63146] = 62;
// bram[63147] = 41;
// bram[63148] = 24;
// bram[63149] = 11;
// bram[63150] = 2;
// bram[63151] = 0;
// bram[63152] = 2;
// bram[63153] = 10;
// bram[63154] = 22;
// bram[63155] = 39;
// bram[63156] = 60;
// bram[63157] = 83;
// bram[63158] = 108;
// bram[63159] = 134;
// bram[63160] = 160;
// bram[63161] = 184;
// bram[63162] = 206;
// bram[63163] = 225;
// bram[63164] = 239;
// bram[63165] = 249;
// bram[63166] = 253;
// bram[63167] = 252;
// bram[63168] = 246;
// bram[63169] = 235;
// bram[63170] = 219;
// bram[63171] = 200;
// bram[63172] = 177;
// bram[63173] = 152;
// bram[63174] = 126;
// bram[63175] = 101;
// bram[63176] = 76;
// bram[63177] = 53;
// bram[63178] = 33;
// bram[63179] = 18;
// bram[63180] = 7;
// bram[63181] = 1;
// bram[63182] = 0;
// bram[63183] = 4;
// bram[63184] = 14;
// bram[63185] = 28;
// bram[63186] = 47;
// bram[63187] = 69;
// bram[63188] = 93;
// bram[63189] = 119;
// bram[63190] = 145;
// bram[63191] = 170;
// bram[63192] = 194;
// bram[63193] = 214;
// bram[63194] = 231;
// bram[63195] = 244;
// bram[63196] = 251;
// bram[63197] = 253;
// bram[63198] = 251;
// bram[63199] = 242;
// bram[63200] = 229;
// bram[63201] = 212;
// bram[63202] = 191;
// bram[63203] = 167;
// bram[63204] = 142;
// bram[63205] = 116;
// bram[63206] = 90;
// bram[63207] = 66;
// bram[63208] = 45;
// bram[63209] = 27;
// bram[63210] = 13;
// bram[63211] = 4;
// bram[63212] = 0;
// bram[63213] = 1;
// bram[63214] = 8;
// bram[63215] = 19;
// bram[63216] = 36;
// bram[63217] = 56;
// bram[63218] = 79;
// bram[63219] = 104;
// bram[63220] = 129;
// bram[63221] = 155;
// bram[63222] = 180;
// bram[63223] = 202;
// bram[63224] = 221;
// bram[63225] = 237;
// bram[63226] = 247;
// bram[63227] = 253;
// bram[63228] = 253;
// bram[63229] = 248;
// bram[63230] = 238;
// bram[63231] = 223;
// bram[63232] = 204;
// bram[63233] = 182;
// bram[63234] = 157;
// bram[63235] = 131;
// bram[63236] = 105;
// bram[63237] = 80;
// bram[63238] = 57;
// bram[63239] = 37;
// bram[63240] = 20;
// bram[63241] = 8;
// bram[63242] = 1;
// bram[63243] = 0;
// bram[63244] = 3;
// bram[63245] = 12;
// bram[63246] = 25;
// bram[63247] = 43;
// bram[63248] = 65;
// bram[63249] = 89;
// bram[63250] = 114;
// bram[63251] = 140;
// bram[63252] = 166;
// bram[63253] = 189;
// bram[63254] = 211;
// bram[63255] = 228;
// bram[63256] = 242;
// bram[63257] = 250;
// bram[63258] = 253;
// bram[63259] = 251;
// bram[63260] = 244;
// bram[63261] = 232;
// bram[63262] = 215;
// bram[63263] = 195;
// bram[63264] = 172;
// bram[63265] = 147;
// bram[63266] = 121;
// bram[63267] = 95;
// bram[63268] = 70;
// bram[63269] = 48;
// bram[63270] = 30;
// bram[63271] = 15;
// bram[63272] = 5;
// bram[63273] = 0;
// bram[63274] = 0;
// bram[63275] = 6;
// bram[63276] = 17;
// bram[63277] = 32;
// bram[63278] = 52;
// bram[63279] = 74;
// bram[63280] = 99;
// bram[63281] = 125;
// bram[63282] = 151;
// bram[63283] = 176;
// bram[63284] = 198;
// bram[63285] = 218;
// bram[63286] = 234;
// bram[63287] = 246;
// bram[63288] = 252;
// bram[63289] = 253;
// bram[63290] = 249;
// bram[63291] = 240;
// bram[63292] = 226;
// bram[63293] = 207;
// bram[63294] = 186;
// bram[63295] = 162;
// bram[63296] = 136;
// bram[63297] = 110;
// bram[63298] = 85;
// bram[63299] = 61;
// bram[63300] = 40;
// bram[63301] = 23;
// bram[63302] = 10;
// bram[63303] = 2;
// bram[63304] = 0;
// bram[63305] = 2;
// bram[63306] = 10;
// bram[63307] = 23;
// bram[63308] = 40;
// bram[63309] = 60;
// bram[63310] = 84;
// bram[63311] = 109;
// bram[63312] = 135;
// bram[63313] = 161;
// bram[63314] = 185;
// bram[63315] = 207;
// bram[63316] = 225;
// bram[63317] = 239;
// bram[63318] = 249;
// bram[63319] = 253;
// bram[63320] = 252;
// bram[63321] = 246;
// bram[63322] = 235;
// bram[63323] = 219;
// bram[63324] = 199;
// bram[63325] = 176;
// bram[63326] = 151;
// bram[63327] = 125;
// bram[63328] = 100;
// bram[63329] = 75;
// bram[63330] = 52;
// bram[63331] = 33;
// bram[63332] = 17;
// bram[63333] = 6;
// bram[63334] = 0;
// bram[63335] = 0;
// bram[63336] = 5;
// bram[63337] = 15;
// bram[63338] = 29;
// bram[63339] = 48;
// bram[63340] = 70;
// bram[63341] = 94;
// bram[63342] = 120;
// bram[63343] = 146;
// bram[63344] = 171;
// bram[63345] = 194;
// bram[63346] = 215;
// bram[63347] = 232;
// bram[63348] = 244;
// bram[63349] = 251;
// bram[63350] = 253;
// bram[63351] = 250;
// bram[63352] = 242;
// bram[63353] = 229;
// bram[63354] = 211;
// bram[63355] = 190;
// bram[63356] = 166;
// bram[63357] = 141;
// bram[63358] = 115;
// bram[63359] = 89;
// bram[63360] = 65;
// bram[63361] = 44;
// bram[63362] = 26;
// bram[63363] = 12;
// bram[63364] = 3;
// bram[63365] = 0;
// bram[63366] = 1;
// bram[63367] = 8;
// bram[63368] = 20;
// bram[63369] = 36;
// bram[63370] = 56;
// bram[63371] = 79;
// bram[63372] = 104;
// bram[63373] = 130;
// bram[63374] = 156;
// bram[63375] = 181;
// bram[63376] = 203;
// bram[63377] = 222;
// bram[63378] = 237;
// bram[63379] = 248;
// bram[63380] = 253;
// bram[63381] = 253;
// bram[63382] = 247;
// bram[63383] = 237;
// bram[63384] = 222;
// bram[63385] = 203;
// bram[63386] = 181;
// bram[63387] = 156;
// bram[63388] = 130;
// bram[63389] = 104;
// bram[63390] = 79;
// bram[63391] = 56;
// bram[63392] = 36;
// bram[63393] = 20;
// bram[63394] = 8;
// bram[63395] = 1;
// bram[63396] = 0;
// bram[63397] = 3;
// bram[63398] = 12;
// bram[63399] = 26;
// bram[63400] = 44;
// bram[63401] = 65;
// bram[63402] = 89;
// bram[63403] = 115;
// bram[63404] = 141;
// bram[63405] = 166;
// bram[63406] = 190;
// bram[63407] = 211;
// bram[63408] = 229;
// bram[63409] = 242;
// bram[63410] = 250;
// bram[63411] = 253;
// bram[63412] = 251;
// bram[63413] = 244;
// bram[63414] = 231;
// bram[63415] = 215;
// bram[63416] = 194;
// bram[63417] = 171;
// bram[63418] = 146;
// bram[63419] = 120;
// bram[63420] = 94;
// bram[63421] = 70;
// bram[63422] = 48;
// bram[63423] = 29;
// bram[63424] = 14;
// bram[63425] = 5;
// bram[63426] = 0;
// bram[63427] = 1;
// bram[63428] = 6;
// bram[63429] = 17;
// bram[63430] = 33;
// bram[63431] = 52;
// bram[63432] = 75;
// bram[63433] = 100;
// bram[63434] = 126;
// bram[63435] = 152;
// bram[63436] = 176;
// bram[63437] = 199;
// bram[63438] = 219;
// bram[63439] = 235;
// bram[63440] = 246;
// bram[63441] = 252;
// bram[63442] = 253;
// bram[63443] = 249;
// bram[63444] = 239;
// bram[63445] = 225;
// bram[63446] = 207;
// bram[63447] = 185;
// bram[63448] = 161;
// bram[63449] = 135;
// bram[63450] = 109;
// bram[63451] = 84;
// bram[63452] = 60;
// bram[63453] = 40;
// bram[63454] = 23;
// bram[63455] = 10;
// bram[63456] = 2;
// bram[63457] = 0;
// bram[63458] = 2;
// bram[63459] = 10;
// bram[63460] = 23;
// bram[63461] = 40;
// bram[63462] = 61;
// bram[63463] = 85;
// bram[63464] = 110;
// bram[63465] = 136;
// bram[63466] = 162;
// bram[63467] = 186;
// bram[63468] = 208;
// bram[63469] = 226;
// bram[63470] = 240;
// bram[63471] = 249;
// bram[63472] = 253;
// bram[63473] = 252;
// bram[63474] = 246;
// bram[63475] = 234;
// bram[63476] = 218;
// bram[63477] = 198;
// bram[63478] = 175;
// bram[63479] = 150;
// bram[63480] = 125;
// bram[63481] = 99;
// bram[63482] = 74;
// bram[63483] = 51;
// bram[63484] = 32;
// bram[63485] = 17;
// bram[63486] = 6;
// bram[63487] = 0;
// bram[63488] = 0;
// bram[63489] = 5;
// bram[63490] = 15;
// bram[63491] = 30;
// bram[63492] = 49;
// bram[63493] = 71;
// bram[63494] = 95;
// bram[63495] = 121;
// bram[63496] = 147;
// bram[63497] = 172;
// bram[63498] = 195;
// bram[63499] = 215;
// bram[63500] = 232;
// bram[63501] = 244;
// bram[63502] = 251;
// bram[63503] = 253;
// bram[63504] = 250;
// bram[63505] = 242;
// bram[63506] = 228;
// bram[63507] = 210;
// bram[63508] = 189;
// bram[63509] = 165;
// bram[63510] = 140;
// bram[63511] = 114;
// bram[63512] = 88;
// bram[63513] = 64;
// bram[63514] = 43;
// bram[63515] = 25;
// bram[63516] = 12;
// bram[63517] = 3;
// bram[63518] = 0;
// bram[63519] = 1;
// bram[63520] = 8;
// bram[63521] = 20;
// bram[63522] = 37;
// bram[63523] = 57;
// bram[63524] = 80;
// bram[63525] = 105;
// bram[63526] = 131;
// bram[63527] = 157;
// bram[63528] = 182;
// bram[63529] = 204;
// bram[63530] = 223;
// bram[63531] = 238;
// bram[63532] = 248;
// bram[63533] = 253;
// bram[63534] = 253;
// bram[63535] = 247;
// bram[63536] = 237;
// bram[63537] = 221;
// bram[63538] = 202;
// bram[63539] = 180;
// bram[63540] = 155;
// bram[63541] = 129;
// bram[63542] = 103;
// bram[63543] = 78;
// bram[63544] = 55;
// bram[63545] = 35;
// bram[63546] = 19;
// bram[63547] = 8;
// bram[63548] = 1;
// bram[63549] = 0;
// bram[63550] = 4;
// bram[63551] = 13;
// bram[63552] = 27;
// bram[63553] = 45;
// bram[63554] = 66;
// bram[63555] = 90;
// bram[63556] = 116;
// bram[63557] = 142;
// bram[63558] = 167;
// bram[63559] = 191;
// bram[63560] = 212;
// bram[63561] = 229;
// bram[63562] = 242;
// bram[63563] = 251;
// bram[63564] = 253;
// bram[63565] = 251;
// bram[63566] = 243;
// bram[63567] = 231;
// bram[63568] = 214;
// bram[63569] = 193;
// bram[63570] = 170;
// bram[63571] = 145;
// bram[63572] = 119;
// bram[63573] = 93;
// bram[63574] = 69;
// bram[63575] = 47;
// bram[63576] = 28;
// bram[63577] = 14;
// bram[63578] = 4;
// bram[63579] = 0;
// bram[63580] = 1;
// bram[63581] = 7;
// bram[63582] = 18;
// bram[63583] = 34;
// bram[63584] = 53;
// bram[63585] = 76;
// bram[63586] = 101;
// bram[63587] = 127;
// bram[63588] = 152;
// bram[63589] = 177;
// bram[63590] = 200;
// bram[63591] = 220;
// bram[63592] = 235;
// bram[63593] = 246;
// bram[63594] = 252;
// bram[63595] = 253;
// bram[63596] = 249;
// bram[63597] = 239;
// bram[63598] = 225;
// bram[63599] = 206;
// bram[63600] = 184;
// bram[63601] = 160;
// bram[63602] = 134;
// bram[63603] = 108;
// bram[63604] = 83;
// bram[63605] = 60;
// bram[63606] = 39;
// bram[63607] = 22;
// bram[63608] = 9;
// bram[63609] = 2;
// bram[63610] = 0;
// bram[63611] = 2;
// bram[63612] = 11;
// bram[63613] = 24;
// bram[63614] = 41;
// bram[63615] = 62;
// bram[63616] = 86;
// bram[63617] = 111;
// bram[63618] = 137;
// bram[63619] = 163;
// bram[63620] = 187;
// bram[63621] = 208;
// bram[63622] = 226;
// bram[63623] = 240;
// bram[63624] = 249;
// bram[63625] = 253;
// bram[63626] = 252;
// bram[63627] = 245;
// bram[63628] = 234;
// bram[63629] = 217;
// bram[63630] = 197;
// bram[63631] = 175;
// bram[63632] = 150;
// bram[63633] = 124;
// bram[63634] = 98;
// bram[63635] = 73;
// bram[63636] = 51;
// bram[63637] = 32;
// bram[63638] = 16;
// bram[63639] = 6;
// bram[63640] = 0;
// bram[63641] = 0;
// bram[63642] = 5;
// bram[63643] = 15;
// bram[63644] = 30;
// bram[63645] = 49;
// bram[63646] = 71;
// bram[63647] = 96;
// bram[63648] = 122;
// bram[63649] = 148;
// bram[63650] = 173;
// bram[63651] = 196;
// bram[63652] = 216;
// bram[63653] = 233;
// bram[63654] = 245;
// bram[63655] = 252;
// bram[63656] = 253;
// bram[63657] = 250;
// bram[63658] = 241;
// bram[63659] = 228;
// bram[63660] = 210;
// bram[63661] = 188;
// bram[63662] = 165;
// bram[63663] = 139;
// bram[63664] = 113;
// bram[63665] = 87;
// bram[63666] = 64;
// bram[63667] = 42;
// bram[63668] = 25;
// bram[63669] = 11;
// bram[63670] = 3;
// bram[63671] = 0;
// bram[63672] = 2;
// bram[63673] = 9;
// bram[63674] = 21;
// bram[63675] = 38;
// bram[63676] = 58;
// bram[63677] = 81;
// bram[63678] = 106;
// bram[63679] = 132;
// bram[63680] = 158;
// bram[63681] = 183;
// bram[63682] = 205;
// bram[63683] = 223;
// bram[63684] = 238;
// bram[63685] = 248;
// bram[63686] = 253;
// bram[63687] = 253;
// bram[63688] = 247;
// bram[63689] = 236;
// bram[63690] = 221;
// bram[63691] = 201;
// bram[63692] = 179;
// bram[63693] = 154;
// bram[63694] = 128;
// bram[63695] = 102;
// bram[63696] = 78;
// bram[63697] = 55;
// bram[63698] = 35;
// bram[63699] = 19;
// bram[63700] = 7;
// bram[63701] = 1;
// bram[63702] = 0;
// bram[63703] = 4;
// bram[63704] = 13;
// bram[63705] = 27;
// bram[63706] = 45;
// bram[63707] = 67;
// bram[63708] = 91;
// bram[63709] = 117;
// bram[63710] = 143;
// bram[63711] = 168;
// bram[63712] = 192;
// bram[63713] = 213;
// bram[63714] = 230;
// bram[63715] = 243;
// bram[63716] = 251;
// bram[63717] = 253;
// bram[63718] = 251;
// bram[63719] = 243;
// bram[63720] = 230;
// bram[63721] = 213;
// bram[63722] = 193;
// bram[63723] = 169;
// bram[63724] = 144;
// bram[63725] = 118;
// bram[63726] = 92;
// bram[63727] = 68;
// bram[63728] = 46;
// bram[63729] = 28;
// bram[63730] = 14;
// bram[63731] = 4;
// bram[63732] = 0;
// bram[63733] = 1;
// bram[63734] = 7;
// bram[63735] = 18;
// bram[63736] = 34;
// bram[63737] = 54;
// bram[63738] = 77;
// bram[63739] = 102;
// bram[63740] = 127;
// bram[63741] = 153;
// bram[63742] = 178;
// bram[63743] = 201;
// bram[63744] = 220;
// bram[63745] = 236;
// bram[63746] = 247;
// bram[63747] = 253;
// bram[63748] = 253;
// bram[63749] = 248;
// bram[63750] = 239;
// bram[63751] = 224;
// bram[63752] = 205;
// bram[63753] = 183;
// bram[63754] = 159;
// bram[63755] = 133;
// bram[63756] = 107;
// bram[63757] = 82;
// bram[63758] = 59;
// bram[63759] = 38;
// bram[63760] = 21;
// bram[63761] = 9;
// bram[63762] = 2;
// bram[63763] = 0;
// bram[63764] = 3;
// bram[63765] = 11;
// bram[63766] = 24;
// bram[63767] = 42;
// bram[63768] = 63;
// bram[63769] = 87;
// bram[63770] = 112;
// bram[63771] = 138;
// bram[63772] = 164;
// bram[63773] = 188;
// bram[63774] = 209;
// bram[63775] = 227;
// bram[63776] = 241;
// bram[63777] = 250;
// bram[63778] = 253;
// bram[63779] = 252;
// bram[63780] = 245;
// bram[63781] = 233;
// bram[63782] = 217;
// bram[63783] = 197;
// bram[63784] = 174;
// bram[63785] = 149;
// bram[63786] = 123;
// bram[63787] = 97;
// bram[63788] = 72;
// bram[63789] = 50;
// bram[63790] = 31;
// bram[63791] = 16;
// bram[63792] = 5;
// bram[63793] = 0;
// bram[63794] = 0;
// bram[63795] = 5;
// bram[63796] = 16;
// bram[63797] = 31;
// bram[63798] = 50;
// bram[63799] = 72;
// bram[63800] = 97;
// bram[63801] = 123;
// bram[63802] = 149;
// bram[63803] = 174;
// bram[63804] = 197;
// bram[63805] = 217;
// bram[63806] = 233;
// bram[63807] = 245;
// bram[63808] = 252;
// bram[63809] = 253;
// bram[63810] = 250;
// bram[63811] = 241;
// bram[63812] = 227;
// bram[63813] = 209;
// bram[63814] = 188;
// bram[63815] = 164;
// bram[63816] = 138;
// bram[63817] = 112;
// bram[63818] = 87;
// bram[63819] = 63;
// bram[63820] = 42;
// bram[63821] = 24;
// bram[63822] = 11;
// bram[63823] = 3;
// bram[63824] = 0;
// bram[63825] = 2;
// bram[63826] = 9;
// bram[63827] = 21;
// bram[63828] = 38;
// bram[63829] = 59;
// bram[63830] = 82;
// bram[63831] = 107;
// bram[63832] = 133;
// bram[63833] = 159;
// bram[63834] = 183;
// bram[63835] = 205;
// bram[63836] = 224;
// bram[63837] = 239;
// bram[63838] = 248;
// bram[63839] = 253;
// bram[63840] = 252;
// bram[63841] = 247;
// bram[63842] = 236;
// bram[63843] = 220;
// bram[63844] = 201;
// bram[63845] = 178;
// bram[63846] = 153;
// bram[63847] = 127;
// bram[63848] = 102;
// bram[63849] = 77;
// bram[63850] = 54;
// bram[63851] = 34;
// bram[63852] = 18;
// bram[63853] = 7;
// bram[63854] = 1;
// bram[63855] = 0;
// bram[63856] = 4;
// bram[63857] = 14;
// bram[63858] = 28;
// bram[63859] = 46;
// bram[63860] = 68;
// bram[63861] = 92;
// bram[63862] = 118;
// bram[63863] = 144;
// bram[63864] = 169;
// bram[63865] = 193;
// bram[63866] = 213;
// bram[63867] = 230;
// bram[63868] = 243;
// bram[63869] = 251;
// bram[63870] = 253;
// bram[63871] = 251;
// bram[63872] = 243;
// bram[63873] = 230;
// bram[63874] = 213;
// bram[63875] = 192;
// bram[63876] = 168;
// bram[63877] = 143;
// bram[63878] = 117;
// bram[63879] = 91;
// bram[63880] = 67;
// bram[63881] = 45;
// bram[63882] = 27;
// bram[63883] = 13;
// bram[63884] = 4;
// bram[63885] = 0;
// bram[63886] = 1;
// bram[63887] = 7;
// bram[63888] = 19;
// bram[63889] = 35;
// bram[63890] = 55;
// bram[63891] = 78;
// bram[63892] = 103;
// bram[63893] = 128;
// bram[63894] = 154;
// bram[63895] = 179;
// bram[63896] = 201;
// bram[63897] = 221;
// bram[63898] = 236;
// bram[63899] = 247;
// bram[63900] = 253;
// bram[63901] = 253;
// bram[63902] = 248;
// bram[63903] = 238;
// bram[63904] = 223;
// bram[63905] = 205;
// bram[63906] = 182;
// bram[63907] = 158;
// bram[63908] = 132;
// bram[63909] = 106;
// bram[63910] = 81;
// bram[63911] = 58;
// bram[63912] = 38;
// bram[63913] = 21;
// bram[63914] = 9;
// bram[63915] = 2;
// bram[63916] = 0;
// bram[63917] = 3;
// bram[63918] = 11;
// bram[63919] = 25;
// bram[63920] = 43;
// bram[63921] = 64;
// bram[63922] = 88;
// bram[63923] = 113;
// bram[63924] = 139;
// bram[63925] = 165;
// bram[63926] = 188;
// bram[63927] = 210;
// bram[63928] = 228;
// bram[63929] = 241;
// bram[63930] = 250;
// bram[63931] = 253;
// bram[63932] = 252;
// bram[63933] = 245;
// bram[63934] = 233;
// bram[63935] = 216;
// bram[63936] = 196;
// bram[63937] = 173;
// bram[63938] = 148;
// bram[63939] = 122;
// bram[63940] = 96;
// bram[63941] = 71;
// bram[63942] = 49;
// bram[63943] = 30;
// bram[63944] = 15;
// bram[63945] = 5;
// bram[63946] = 0;
// bram[63947] = 0;
// bram[63948] = 6;
// bram[63949] = 16;
// bram[63950] = 32;
// bram[63951] = 51;
// bram[63952] = 73;
// bram[63953] = 98;
// bram[63954] = 124;
// bram[63955] = 150;
// bram[63956] = 175;
// bram[63957] = 198;
// bram[63958] = 217;
// bram[63959] = 234;
// bram[63960] = 245;
// bram[63961] = 252;
// bram[63962] = 253;
// bram[63963] = 249;
// bram[63964] = 240;
// bram[63965] = 226;
// bram[63966] = 208;
// bram[63967] = 187;
// bram[63968] = 163;
// bram[63969] = 137;
// bram[63970] = 111;
// bram[63971] = 86;
// bram[63972] = 62;
// bram[63973] = 41;
// bram[63974] = 24;
// bram[63975] = 11;
// bram[63976] = 2;
// bram[63977] = 0;
// bram[63978] = 2;
// bram[63979] = 9;
// bram[63980] = 22;
// bram[63981] = 39;
// bram[63982] = 60;
// bram[63983] = 83;
// bram[63984] = 108;
// bram[63985] = 134;
// bram[63986] = 160;
// bram[63987] = 184;
// bram[63988] = 206;
// bram[63989] = 225;
// bram[63990] = 239;
// bram[63991] = 249;
// bram[63992] = 253;
// bram[63993] = 252;
// bram[63994] = 246;
// bram[63995] = 235;
// bram[63996] = 219;
// bram[63997] = 200;
// bram[63998] = 177;
// bram[63999] = 152;
    // end
    // // Initial block to load BRAM (use this for simulation or pre-synthesis testing)
    initial begin
        $readmemh("input.mem", bram);  // Replace "input.mem" with your file name
    end

    // vars
    logic[31:0] f0;

    logic [7:0] audio_sample;
    logic [10:0] audio_sample_counter;
    logic [63:0] audio_addr;
    logic audio_sample_valid;

    logic start_computation;
    logic f_out_valid;

    logic [6:0] note_num;
    logic [5:0] band_counter; // waits until the audio sample has been run through bandpass to send another one

    typedef enum {IDLE, LOAD, YIN, UPDATE} states;
    states state;

    logic go_update;



    // audio_processing audio_processor (
    //     .clk_in(clk_in),
    //     .rst_in(rst_in),
    //     .audio_in(audio_sample),
    //     .audio_in_valid(audio_sample_valid),
    //     .start_computation(start_computation),
    //     .f_out(f0),
    //     .f_out_valid(f_out_valid)
    // );

    yinner_song audio_processor (
        .clk_in(clk_in),
        .rst_in(rst_in),
        .sig_in({1'b0, audio_sample}),
        .sig_in_valid(audio_sample_valid),
        .start_computation(start_computation),
        .f_out(),
        .f0(f0),

        .f_out_valid(f_out_valid)
    );
    
    // Read BRAM and store results
    always_ff @(posedge clk_in) begin
        if (rst_in) begin
            audio_sample <= 0;
            audio_sample_valid <= 0;
            audio_addr <= 0;
            audio_sample_counter <= 0;


            start_computation <= 0;
            note_num <= 0;
            band_counter <= 0;

            state <= IDLE;

            for (int i = 0; i < 31; i++) begin
                results[i] <= 0;
            end

            done <= 0;
            go_update <= 0;

        end else begin

            case(state)
                IDLE: begin
                    if (start) begin
                        state <= LOAD;
                        note_num <= 0;
                        audio_addr <= 4000; // change to location of first note
                        audio_sample_counter <= 0;
                        band_counter <= 0;
                    end
                end

                LOAD: begin
                    if (band_counter == 0) begin
                        audio_sample <= bram[audio_addr];
                        audio_sample_valid <= 1;
                        band_counter <= band_counter + 1;
                    end else if (band_counter == 10) begin // arbitrary
                        band_counter <= 0;
                        audio_sample_counter <= audio_sample_counter + 1;
                        audio_addr <= audio_addr + 1;

                        // if we've hit the last sample
                        if (audio_sample_counter == 499) begin
                            state <=  YIN;
                            start_computation <= 1;
                            audio_addr <= audio_addr - 499;
                        end
                    end else begin
                        audio_sample_valid <= 0;
                        band_counter <= band_counter + 1;
                    end
                end

                YIN: begin
                    start_computation <= 0;
                    if (f_out_valid == 1) begin
                        go_update <= 1;
                    end

                    if(go_update) begin
                        state <= UPDATE;
                        go_update <= 0;
                    end
                end

                UPDATE: begin
                    // need to update to next note 
                    if (note_num == 8) begin
                        state <= IDLE;
                        done <= 1;
                    end else begin
                        note_num <= note_num + 1;
                        audio_sample_counter <= 0;
                        band_counter <= 0;
                        audio_addr <= audio_addr + 8000;
                        state <= LOAD;
                    end

                    // and fill the frequency bram
                    results[note_num] <= f0;

                end
            endcase
            
        end
    end
endmodule
